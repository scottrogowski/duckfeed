��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C����FQTX5��)w�"��c��Lg+Z�fvV@4�ZP�>l���
�U��������tAĪj�k��V����>lv�C�/8��M�jR0�:q����Tԅg%�L�:�����t}W�/vF�XȰu���*_=�Ҧ�/W �W�J��k2|�v����Q�o�2�l� �@��n�S&E����q;�Ǹ�(�b�?��&�pAM�� k;Eb���7��U�U�k�и}8�+9$��'����ݧa#{�~P�C@�u`�#����]�S�N{"C=l
�i��+*<�L�n�k��STA��s�%�X;�y��@����L����n��e���-�4���=���t�X�	���B�`�K�C���Ɍb��8!5te���i� �������9�E�y�w��ܺZz�
�5�_�w�.W%x���|�	
�Z�� /��x���f�-H>��|�)O�(�x��:E��&��Ͳ�Q����<>�E������B����
\�t΍��9��Ȟ��\���$�z`�� �1n@4/��e�P��$���u-��?�J�$?���Q�Mʕ��[��y��ن@0ha,��t�H���OD0�p�{O��M=f~-�G����(*��!m�Es'�#�A~�G���yk"�ї�����!A.���Qձ�&Yeis?ޖ`r4��9��7H�͚J9i�Ň�yʣ]��,�y��)�Wz1����?����Wt����� ���� �mT��"�\<��o�����D���^ϝe�x鞾�F̂���ˁ��ͪ΢:yz���Jc
��CN�!=�,�]$a�����Ù���2���rTc���Z�=HZ�$�Z��^T�{)�ȧ���_ׇ߹k ݧ �dظ�z����*����D��٥=ɬWb�	օ�����^���Ar�pLPH�7��G(�.O�]\��Snf�ǯy��(za:e�^������.�Ƭ�r}�GMP�s �Ǭ�����O�x����Y�T��3��`��3h�s:����\2�d�;n-�q8���FW��>3�|o�
|�ÿ��F4I����[Lb�8��9'�Yj�l���[T��i�V��p���eƤ��h�9���`=����[Pf��c���#����4�7����Y.@�ݧ��{��Q�MDm��D������C��2��]�4���vK��B����s�6'.s;�Z�U�e9J�:9�7��@T�_��ꐜ�M�x��>�`�� ���"�k�(V�я�����5��GS����ׂk�M���I	ǳS��Q�N��P�ĜF�GA���Wy�j-���D�k�*��M����ՒJ	�q���Y۩>q�S���R�(Em�F��\���-�h���Pj	M4oı����DN�����(,�,�|��SO!A�5��.��2�ɉz�	�K���q�'�=[ʭ|LX��Q�h;vn�S;̝�Є�%/o�f?*���[�B*�z��K4��)�D�gz��+.ݕ��c��%�V{X,,7+M�0cc��;L�W���zo��ϖQ���"�L7�k��1�鲾ě@�uo#]��` �00�v�3)��e�o�g9Д�(�e�$��5�z�m�7*'��
�.�J��ly�L:,ۨWu0B٤����?��RĘB+%yY�|�Q@������¯C>�<卓���<X�dI���I:�!�r�4+#(lpؒ&1���эb_�+V"������a!!�h4�B��PS@ {4�i.����eG�\�w9v��<��pp풥�OYY�0������Co�gFFp�[�|o�s��u��-W/�Hx�o3p�+F�;Lг6]6b��$�^W(�,ބ$���(�?�g&kyt_�e���s5���VE����{l8ݎ��Z�x�'8�^+��Wl8˧N�]v�Xѡ�t �m\K ���a����)\�$J{�[�=�4��h�}�iy2Z��TDy2@��k�N0��~���qt�x)�{��N<��LW`��uT�*���(�;�)��)���@N{��'zoT)G� B|e�eH\�(8���@�,�V�6����r��_8K�E:��&w �aeC�&f.f\*������2�e��C����<���
0�?��u\kYA^M��*��i^�X	��0]Zs��))�z	��l��8k�aNe2��i��3V5��]��zv��� f�\��$��Oƺ����Ni.�q-�Ӭ#��X�	O6�<�)��c�Xͱ�3��X�Qw���8RJ�x�(��xsC�-�
;Տ����px��'lHR
��Z��{|�{�1,
 �e7ų��	f��������~�GPV�S5U��0���(�ẗx4��������W��H;�*����j�;��������f�������D�Q�H�Nڡ��gT�Aw75��7�:�C�X��4�>�<%�i�Z;n5�VJU}!�0��zu3���ky��`0��M��
��j����eqw��T�xvB�c�1EzhMP]0X�X
"4p@HHW$�ik\9��D�{����i��Ԉ<�2M�v���,�@-q�%v2���,�=��埱�lѕ#��
%Z˓u��O�
�q�:0m����K�Pu�!0�;���j�\�Kyv�k[�0z�GN����ժ��R�Y8-&����i�]d���� ǹҷ��c�&�qO�&o.F�Eg�=A#%0`�Jn��U5�I!�d�l�J�J���V2Ylie�K��:_BĘ���;�����.B�|d��`�g�- {�y�Jl��L��&r�6 x�M"�p{�[�{Wc�=�!�ٓ.ۓۋ_��I[n^�� L^�
��2���I�R@쒬���H�n}��ఉ�y�fÅ	���>�,r�-�-^�<1�L��$��h˰���L��X�ibI/�K�J��jXc�n��w<�A�J��ȅ?����N�ݤ�z��5H���ߺ�=x��S�ˉVH�x���Ր����p��O(#	�ӽݸ�� '���⩊<0�v�o����V*��Kr-�I
�w		Ŗ��i��|����9|��N�3�
(=��0Sh�@˔��f��Un�6�V5Վx����o��B<�99?P.��/ H����gY#0�<	��� ��+PZ�E�V��)�J
��s���.�N�ΙyŽV���_I��O,��`�'��<|��YЗ�[�QҨZe�T��B�0\�R�:�&�>�B�Nݠ�,ʝ����/��� u�=A����#��d�
z�U�x�5����T��4�sK���m��E5�rfcg9bx���ʶN��V!�Y������)#-D�+)��9D�$���+iV�9�SaP�	�p�~>r�o���n17�7RRZA77e�)*D���˄ߣ�d�f��������)�%��< J�v��)4nO�D�Q�)�wDX5�@a��=�;�7��a_w�OR�zw�r睟�;1�?���17�0F4OaQ���܎��Fk��bp�k��o{��u�������?z��dl�+�H[m��5��xg�#3&4}����J4�
(U��Q�-���3x�T&4H��(����|"��Z.��
���hN���Llk~n�q�A��1��x��Gޓ����bt$���pԸ�P��K4Ķp����w�Kf,8{k�dA�i�p7��֩�i�~}�G�d�Jn/��1?>�n,�i~�n�sh��D���g)O5X��u$+�f���V�z���\(xL՝\�GaIrE/`;�&���m.�7
�\��y4�Ie^S��/u���V1���?���B�e[ '��{��SB� *6���k��� KR����z�����h��g�x�ǭ�ʧ�Č����J;)s'W=w���z�9Ich)=�_�#8�{���\����=�/�`/����ԂapQ�����X�+�^j���`0H�t^͋�Z���u�R�Nl)$�^�w�*<�xG����.����Y���Qp�wu�y`����R�Zj��@�ery���y��	ܠ���w���$�]u`1�f���pd]ӏj��u��&�fU��¤��7��K�>^FA@gp�
��J��N�l��[P��k�Q�����Fy���Un#g	��g��'�mO*��P���N���1�>W��c��l����Nֈ�=��k���6�fsm;�\o��m$hjAW~$��a��o��`�@�c�=7»9u�{^��%�ؤv�F|{c�;ǉ+ac B�f�R�3�g�S��J�Z8�)р���F�OA'y�[��⫖%
�L �0�}żА�f���,^���kи�>l���Hf����j��G%�=�ܣr����dYD}q �y��Hf�
x����F���8#�B�R����s�[�m�Ow�C��"���F)�ޜ6iP��k��ӹ�z����T�;�o�Q���×HE���n� ���z�f��?:N�s��(�j��W*s��u�f8}�U�K5�#a�5+��V�bKI�R�K�rQ�a|�U]��xq�����n���]&%�\�/�a^�:�3Jkc�'l�n��ǎ�5(0Hש-�u��J�z{���@�1Wӆ�̀��������VCQ	K%kl�b.�<�Sx����c�Ü�B�w�1ڙb;u��Ʊ�������50X�hr2�G:�����JI�'�IO�V;Q)+�V���.��wh��.4*�gH:	�(7-��[X�DT�L���j,ӏ[���e8�'xd�O���*���Yrnx(������x&,K�<���d�SU�ߗ��J	�7��J?H�ڒ�@�f�p�"ћT�#%�E/}�K����>:E�����k�R.��Q/��7���%�ʪ�b��|�/1�b���谕�TS���~���*�5GKf�/qk����F��TkF'��ReY�KmVv/����-B2 �`��j$����M�FGC�`Y����EB�I�e����P]N/:��9�_�����N.��s��s���4]�aI�5�
�l��N�M��5����W�!�]f[���h1Ħ	��Ń�_ZX�l�է賁�U^Y�E2|��lƉ��^[)�G�����8�%2�0X�D�t��¿?B�O�7���ū̠�8�N�"8�;-�j!����Wk�}/����ȳr�6�(�e�}T��2�U�P+@ސ�ӆ���AϮ�R7D�D�/+��oC�1�U�#�i��_p�4�3��G%�]#��NwN�zY��Vۧth���������TL�`�3g�;�e�a�@L?���t�mOWX�p�s:�V����a�����C�!_�I�w�)���a�������xُ�+����R ��(T�ierUc�4���t+!��cO0=n��+�CDp�!}g0��I���jH �A;:.4bYv��#�w�O���c9�@	�K�5���Z��
�$.��c�+���cr�3d��$Ч��ˬ$�G�-��n�%L������Fdi2������t�H�y�,���v �$�=Ͻ���9��[��r��5��9�J>��T,��X����ʟ��EQ��)|,��C�]8�����y|dާ*��D~����#Un+~.�$�x#b��v4����v�=�Ohيr_���1敾W�	������p��1�t�.4æ�e4~��"8/V������|*������贼�((@��]{Z��H�� ���\�s�w�G���q't����[!`t,wNV�8㾽�-_q3��hD�6H���%fv-��4���a8��5�N:�)�[���_l��F�yXX�������+��x&`,��Z�`��7?g�/b�ɀ �9����/���o.1Ʒv4k=��z����Xn���0�Y�4!���A�!���mK�{��FE��Ww8��qeVd(�%J¹���0��ܹ��;L#0ݱ=���]P�j��"]��i�CC�&�GZ�VY�+#C�a�@E@���2�� -"'�xf��s��6�mY2.	��P/�G��$s|��AU.�M=��+p«3TF�Y�@t,�Qb
��5�Xj|�*8��n4�]��ii�l��Y6,c��1\���&�����k���e1�m�<������T�=:�#��Uy:2�� a�C6�0�gܛ�q,Ix����Z����-�e�JB� jnJ`��~�1�q��ڀ���2�j�Q:�@?b��1��;��,x&b '�8?�`S#��B����&��iB�]@�L�#�/o[�oI�
�:�4��o�ͬ)�K���@��
Nf<$���m/!�"�׏��3� �����T��Ƒ��=��y�-�r�1! ��1ix_����v�3BR7���I�]��)PS�ҧ��f_kA����Q?m�������hc���P�z%��,~k���w�Ͷ��Ξa�Q��ܪr/�t�EuP���6�f�������a�����W_�J@KL�9�`�#��-疩/bl�FW!1�����*�����wZ�)��f���ԃ��J�A�.�h�@C'�����*�T�~��"=��rL' �vC���I�{�- ���&!K(�.�s�����P-��4�Fo���E��w�s� ⢽]���-\O'�߹d�U�	�jH��ԝf4�;rG*D�_6������~P!Z?�;wА�T�T8]�_�>�)M�����tXz=�{���4��rץ(i]�v��Lhϟ�fś!Y�K��m#�/���~�J�	����*�o#\�H�!>3}-����Nl��M�m�__o�`���R�5���R�e���'5Q�Yo����Ø��ԡH��U��t2�o�	�		�*��c�lxe �WEmK��z2��347Ԛi���䩰��bl�Y~��f��Wؾs�ڝ�&Ϳ�	���~'k�gC'���&7K� ���œ9!�;�Ш�"�9����SrEƷ�������Wo0�f%l"�A�M������Nx�9�~#�-Oy�e������Yʛ�=P�[\�o���)ga.�� C��߶gk	w\���w9~l��z5Y�ڻ(�`��,�U����<����kd<"�Fk����i 2�*߻�����m�i����*`��Zɕ��:+�5R/�,M�lb�O��.�� �s��ۓ�e���sY�j�w�P�ku�bm�D|�G'���I�;{���n��&�&��{��4fk+�[���0#��u��%�YǷ���D���ޜꤲ\yjK��~Ɯ��1l���
������i49��\odf��'����$�ۤH;�R���}	]G���T��uZZ�{@ߒOzQ�TY����!�z����ī�jL�n��m����4�sEu�Q�-�	�,5ёZ��C�*uɇ��?'�G�;Ek���ʣ�[��f�;l*�д�#�斡�{��߂��=���"�z��KR��r8]��D7X(�ﴥ��"K��$��|Ao&��v�����75jV,Nh\dΞ�� �I�%h-��C���Yy�1q*j���qN��~������]gG�L�m"k>�����:\���٦' �O\����E���׊���;��;^&ժ�k�P@�·3�z�eȲ-�N \�|�}"�h�e0�����'M�`�x�R�U�"��6�ܳ��ou�ȋ%C��������I�<R��������N�@��J�ٶ�٬�u>;����x��ýCۦ�25�N�S6� �dS�b�y������c���U>Y[|����W�D�;c)f���YY��ELtN]�wg]���.T�c }�f��$tեn�����Y?W�NO��8�w+~]_�*���2�x�e�bq���F��	��bp�$��=5-譖I-3��Bj�?"!�v���A�Q��	��%��c{>o��!�Vޤ����j����b`�P�w}� �dJs)׍Ci�Ej��$��wk���\�
����.8ɲTݑ�^�h��L��?�F��a.dZZ�d�f'gF�7d^ h�ۈ0�I�汓�=�|��^kla+�O���N
�+�S�>zxM��d��U�P��{C�L�Bv�v4̿����q���\��k�G\)/ Q砷D�ǌ}��I���1�&�����ZtN�*�H>d	�3l�V�@��`]����Q��YU��1�#K��?N&�=5��|��ž�%1&���u�)�T�ڞ��p}8��o�����y#�)�����5�5:�'�ũQי&�'��5h��{ֈ��|Q��8
�i �'Om��CK�w��=Vlos�n���a4H&+ؕ�n�{g�|VW�W���LÌ\�Ne%΄�X��h/b-�k	�joz�.�Sn�k��!Ƭ��6���Z����5�;��x@�~Q�˙�ɿ%��='�3�{#���{jᚱ���r�f`��_��+5�&Q����� +M�/���g�@�񡰧�Q�̽U��ꜿC���;��T]�a%S����y�e�e����5:	����b�m�.��Z�5�;;�a��EZE�o�N� iީt�������V^7d�pr���Rʉ5�R����W�5C	�R�y�y<(�wH�o?����.�Qp�DK�}&HG��38\h��/o�\��w<h���Dd;_�cїlX��D�^$/�ۭ̐ߠ��E��?��j�Yz��OE¡՟!U��@S}�G4zj�m=tr��0����ۼ H
�hՄ�OZM��B+���S�(��<��E��>�J�5D�k�0otN�T��Q��Gh�6���^ѷ����3��p#j/�O���� 7���n؈QXܢ���w�u��c�AX�^O~��'^�I3h]�����4sώL!Vr�7��	�g<8a���$i;�
�{0�p*�}�vv��#q�9y}֎6b���l'�Ә�D�Y�EfX�@������5p�����s~�������c�?�4��Y����?��*�s�PK2 �x���x���w��)���X��\��f��K��""�Cx���y�$~�BRvݧY������*�xUhnrY*��Z�U!�%X{�
��T�F�H^툉��s�
ncX�춼�7��\��w�v��$�T�)��w����yp����ICXuu��H�f�:�ִ���<�*Ӭ����9���
���B�ž _�ݥ����HH(C^�#-;��KZ�%�ǐ�D>���?���-9�9<Ԥ��u����_��E�[ꇘa5/Ia�f ����"z^��}H�`첒-�k�)�u:٬9�8U�6�ݎ�~A�E���D��z�h���S��b�W���A��n����*A�%�sf^ �2+�{�by��uַ�#xt�~���*� eT����N�d�����ms��+c���
[�*q�s�*��d,�b�M����͕��7�h���e���{=#�����]��0�I�q8n��h<�P����Q�O���,@4/lS�PZ�ar�&����ƕ�X�=��-P<����&�c^��d��;�`��Ve�^�5����'"'؅�X)(S&�z���J��<�vT��`�'�q�Q�a��%��6Ϳx0��hȡ�pO *u�-��Q��	?C����u����E�C���O{R>�;�Vo��]�J�~��5�:f~. ��r��ͥ|s��9T#A�g����.�����~r������96�7SROT��R��g ��KԞw���G7ߣ�6�u�tn:&��6��|l����K"�(�&�|� K�'���{|f���-ؚWy!��8��?۹�K�\�U���b	��v
�l�������WWh���x�H�����es��b���#!{%����*�-}�{NwK��RۿiX/�Z͜p1�o��nma��-0���;+��t�a�j��4Մ��i4�i��X�rp"���W����S��d椗���%�?�g/�9�c�p��x�4�w
�7@Gpr�P������o��epvRK���J��Ҥ?r����''x+s	|m��;�v���> ���IYH겆���6k���L�O���3 �^a�%y��P��+;��u��yg�`��+k\�������p�=*y�j��r�
��C#�<�^r����V�dv�r��X����!����сj-�[���.�./��T���;^����/A���0�r����3����q#��e+��V��E�L��~� ��h���}��H�]{&k>*��l0�Ne#�b�)�ҕ�8	A]�{썌��*�ʠ<�.K�fVe�fS��*63�5Ӟy�4��?�R�9ǟj�1��_���Cb ���PF4��@T8�e�����1߲H��W��gY{���)�����і+ח�lgk2�������6wq���)��v.����Y��Q� �>	�&q�`�����S������g�e��&����&6^ོ���ir�.(����r6uJbF��\oGo�
�bE1P��/�;M��6-a|�A��T�('Q!
�T�v-�S!�̈́_�9��b9->oM|c"�Y\Tn����df��+�*����-�:ni��jM�7座_��B�^�u"ͩ ��%4�s�I�s�z������z��c[�4��˦��7����+�`���S���#g�~�`�@:�s1�g2�p���[���k�$�V�ɲ+x<h&�#��fp2�A�A�7]����Y�W/%G�I�1W
��\�s.�Tu�t~kdW��~�-����Mh����=ܟl��QV�51�SX�,�]�fHWU9�h���oa�՚ ���
J��t�!�;H��~}i7�<�t�0c%D�>��q&;x�F�d�f�n�
�w�Iȯ��i7D�R� 3�p&�%��F�m>�E+n��FI�eϒ��GT�8F]?�e���rV�"�6I�W'ĉ�&dMP�B�5���5��:~��A�=j�2F�(Ø-�կ�?�|e�#2��W�nE���I���C���Q,�oe�շ�)b�!B^�h�km���L���(>���Nk��ۉ�b�Z�/e�TE2�Ͳe��6`dv8��k�����Q��j��Ks�E��q�W�Uc�"�XYz�w%%#쬏6Tx�����
���L�� $��>�;�ѻ�������ϧoe*���S�"�ǩ�E��y�8$
P7!,�E�����
�!+�Q9�c�*�@o�D�L�߫Q�Es�M���<�n��7�F�t��A0kI�Pg5����0!ͦp~i1�lՉ��C� !w< �� �}�����o���v�ҏC(;������`4wϪ^��An��m0�� �=?:1���e�-�9�mՄ�CL��g�e9�>Bv/82,�xgS	���@ ��Ly�,�����;�L'bzϦn!�g�wG^�f,c�N�/��	��N<@�k�.s�\���B�~�7�)c�GM6J�qW�]j޽�Y��Vn�ږη=yL����o�]�S6ĺX��c/a���(��.�t]т�_P�G�<c]��/�L� ?�����"���N�upwMٔ+	��fD��N��e�L˥m.��`�9Z�۰C42�_
J��B/��v�XU��L����^r�uv�r֪�-Z��v4����)r�ۣ�:4�����?\��eD�6"�4�̠-�����!V�Ug��y�9r�ujpXϽ��a�sP.h�JS��T�]��B��v�r�.ѕ?��m�'O��j�S9̌v���4������6�X�8׌��H�"p6yYF�q<�����Oׄ+��nZo��h�!�[.��b�E����`E��K6��n(N�n튱���2�P���c�'��������V n�
�]>�e��˓����O���fP�nN�Vgc���w���h�QBm�W�N��T�Z�wCX�����W�#I��W�Z�i���^�,.W��(A�C�*A�,#�>aϵa!�L>ۅG;f�=+*(����]����ϫRV�Ƭ�Ǟq{�gY�������<! d���+3�>��[�)m?��N��z�QLZ[[(M��w�ʱ�\�6�b"�޹|1Ȼ���FV���T�DID�p$+aoc�P:�t͉n�����a� 2�G�ż�����O9�=��I���T�1�S�Žp���rZ�0Q��NK7�2���N��vD�ێ�z��$2z�T�F�b��@�@o�;�I]��y���=�3�_������yd~;"�<����Y��P z�b��8Y��l7>���ϧ{�(+�q�Y/~Xt����$�.��{Ǌ۲F��m�4%Ѯ�����*	@U�"���?j֞Y�+V;|��VH���T���d*���S~k����_>��������#e�	wC_1�&�ў�!���~͹���[�k��2h��{h�UwW�>|:0�nȈ�FGe͒�%��'�����e|����b�]F7�Np,r����5Fd�!2|?�����`�i>VMT��X1)E�������p�c��*��\rfݽ�c�QsmY��J6	�q�׋V�fK%r���h��ћ���ޣI;�b@A�S+�Rqb����o_"C�������W�J�/����59t��Gd������b�<&�9�ߤ�$�N��5Z}�����U���W1�ӽ.~�3
?t"���H����T�s|��Y6�d�����N�q���bN����D��ŖL%��b���>�T�ٽ�4%<C�>W��f��`s#^���@I��dl-|�׼��0��&��K=*�G�C�kX��T2�k�RMI��Z|�����ݍ�j����6T3�����^f�p� ����~�U���:7;�f�S'ep��^�N�D�Bs�����k��%d�laB��O���*�����x㚶�wbj~�G7a���� ��)I�?,?3р�%U(M���%��6��!$e�"�:sUX;^2=�x�h��frș�����>	e�~]�U�1���\�:�2R���A;]�%�*o��:���N��Zy�T�����`�=?���Sq��JW�O		{�- w/#�S�H�P��/C����?R3|���й�zmO[똿dkfS�!�޳<g�V�a����t�N�V-� �eȪX%b�(�)#DoN}T�xNW��52Ӭ�܉�J�-���3��'���r]�DyGC&�����n��Hk�9O�[��#�����̣�%�w�C�+x�pi>S�ȑ����������~�'��+��Cv�m��IX�)n��R�"����Ƶ�S���)]G����[����IF��Ѿ
L̺�Ke�J��,�i�APV������K����a����D}h����S0EAKTCK�]��j��?�sd��A<C	åCW���NE��6	aΛ���./>��k񊯚p���&�?G�sO!,>W{��v��w=��ZJSz!*3��1*��Q���҃�0�ڐQ��m�Hΐ�3-�Mx��\�G�eQy~��#X�4ϟV��%YH�7a�0�7P�\`Q?��5V<E�*�xН��r�Z��[9nv��Z�Fb���e��8�hd�����+;:P��	�'�O����J/�e����ޮP��w�t>��k��	�����=��ɞ�*��H;`��Ǹ�*J���b�*0ko�7�W0^քىSKVzה+n�����F��tk�wh�e)Δ�m��ʝ
�Vv�k	�����
R�*3\<jm�P �pX�l��m�bڪ��J��^��������6wq��:"�TQ��(k��A�m�VlD�o�7g9�Ri.kD�����Q HdP�/p�Gw�PXTEB�&��/�dGCn�������u
�63��T��� �����{�f !;t���g������R�8�6�a��k����]��ܭѴN2�gt�6A?��YK-�$���@^}<��m9(��#�����cy!$o5:DC�ev�B����F0�'�s�1HG�	1o���Г�X����r��>��.�IPY���5�� ΃�8�\�A
��0:������_mbE�nM?C�J
����Dm��e7sAs��s�sfR]�!���F/�C�8�ܻ��)ҝ�?�s[C��x��TvBN�+.�J�ǋ��n��nkK;L,,�{L�i�i\}pB�T�B�S�}���-�M�*����0��#:�j˕! @��Me@�	9w3��`�a��ޯ���B#ߴoҵ�b~������Z� F,�ŅҾ��Ē����q��kJ���_�)��Vv�ת?
_t=�2t�1OoH��'(+l��^��`+��7��RΈ�0��7&U�o_?��'?�v�0���\O�!�<raa����n��"�_8�c�Ժ�u%~;��Q���kD��K�%V��E��^��_�W-��:lUđ���3,T{�V�Ou^/YK�x�gD��d��"3�HMkX�?�|��äje�=��;9��;��h#�f4���k�u(e���h����g�ȍ~�����e����᳸�hS�0�L�Ӵ
�R_��PE�b4�C{�99�ky*ɮ3��*���±�K���7�G�dv6��>��ہ�l�'�_cҌ�� 60��ZR�@n�j�m���꼙9+�5�*��E�h�'.�CC�6��f�|1�Ǒسp�oȬOL�N����.%�Fn�j�=cs����[���S܇��S��
��v����|��o:4i�
�X�<g],�{)�G�!��g�uV�3�ѩk���ٍ���D��]j���ғ
xL��;#�i}NxR߳��*5:I�Ȫ���� n1��gy�7��FW�tԩ�AՁ�wh�ěҬ� �"\k��#o��]���"��UP�3a]�,�ү�}@�I��RJ<�#�1����� ����դ�@o1#߻����ܠ�h}�o���3>�r�ks<�G�r��<�@�	#���
�����D�J�򘩴h�6��'��ȏ�sе��_Ri��%c�(��K�O"*AR3ϕ���)1�L z��l��~�Fu?���@Y I��<ʄ�a�'�͐����1@�|;���gw}�����X�7��)��1�9|�u\���-�4�^���	�A��]��m���l\�Nc�A�Ãg���uk��8⿈=��>�� �ܟ!EM���j����K�,��ߕ��"�,4��3�o, 3k���b諽sN�E~$6���>�b{��lɞ�����`��Z,���gB%�&lX���� ���E.��覸�ߘ_�e?&�]�� E�pS�˿Q#䔬���WUX!]�v���LIw&�,�7�u����ͯzU��6��Ȓ�[�'REd�\5Д�dϨH�H��, d7Rf�>�c�7�<o�\$<0ܪ���_9�h�q�IA�Y��*��o�l��eB�M�?̅���c4�D��PE��x�tDA����W��H�[D�ޥ���Q�>����\n8�z�!}���@�#n(�N�N�������\�ך���<���%���3��?m]�QM1bW�����d���xL��vnYs���;�n�:����,�P��TZ�e!��#�;t
��꤭��vf;� �=e+�&N��ߺ��QY�D:��-�p8v|I��N��˭�7i^ݱ>Vf���j���,�E�u��� {�N���pOVb:�2���czhl|��YpE��+�DG�����3��[#����*5�f�'�fl�d��YZ<ȧ�z�͸��q�3k���mg��!��!NC��/��9�����F�>w��Yғ9�={�l��,���Q��Ϛ���wޓҭgDP�����1�����V�1M-0��^�e��/�:�HZ��beQ#�(���ǧ�Π�i���f��垣��	�P{�B���9�('�"O@9qX��7�� �W�,�M� ����g5�I��r��Y������٤x�P�[��
&�h���ә�bU���;���HoHg�į(�W�c�#����`1�{�� �r�̺D#9{��<������"����Z&���r�>	����M<a��}}7xh.C����b[;k���3釮�mԓ��aL҅����ԯ%\������n�9v�F$9�56�n�dY�sq_SCOw�UY��?� ��T>��\����F�����tE�|������a��N}�}i��&3�Oz��AY7A�Ӕ�/���f~�&����2��N-�H;�(��IÙ�!t��Uؓ�{M���hM����e����ʙJ<�m����3;�H��
R�+̇
��??�̵?�ߒ�/��n�:]�9��h�� �O�p�l�V���E��^�]�mʨc#��+1j6p���S�"|G8#jf#�ԄD�R�F��x��d�;�ɭ����v5+�z����Nk���fZ-۶��H�6�O�J����V��[Ja�q��3��e��_�����"� �[�:��|��?D�D�[���=��|��:�0G],�B�t���n��M��v~̮��G`WnHY�i��О'\g?�! )ίR�k |㑶ё�9��<E����?��Or� 0�T~y ���i�Y�R/dy<Z����j�{U`(�W)ǴGv�RW~�ǅ"�Ѣ�*����R�e��n���M���^�Fo\7X����y���KN��Д�Z�
L.�7�a���ڟ4 O��G\
��{��7,�u��	z^S���O��I/�w)[���5�sZR���c�̚�C9ק�ք���ҡI4!��!��D��7�Ɂ����-�2�]䶙��Ə>�~)f���KU����8�[-�ЃY��� ��������$����f�W�8�p���m<_�G�[7�A��P{O.|�~��#��ik�����bʨ��Z��T���N-ՃJ��U���@�CV�-�mP����yU���$���,A�Cl���yd&�'L��=^�Z���ħ�G&.h�	4�ۍ݌{��z��0�f����*գ#	�>��c�sP��
O�s�F�����R�s�����ܡK���b��!��r1�D@�L^ɔ�7k?�#�N-��|܉��]���(ғ42�y�T".�;�"E:���3���܂yŃ�ό�Rۆ��s^�}���3T��
�uG�����_~�p0�n*�ɔ��pl�K�R���`�H �gT�����	@���*E ܇���2��{"s:��~�}V��?6�u�AKW�{@���Xv�7
AivEQ"��B��T������I�I��]'+a	�L#����U3c��Nd�|?Aw*�E_�o��F�A(]7�GY�#��]���U�:�v��.K�d�1�@G�ԥ�9~���H�G����]f�T��r�O�3���O�����%{BU��ղq.�&K	��v3c��\Rw�fH��b�e��Z0v,�l��G cP�K��N���<��:z��
�Fj�!�r�(
��;p�S��D���x����k/��fn��8���5��\��Mv�_e��sF��\SM�r�X���1j�k������*���=�N�,B>�:�5�欏��1��Ep��۠y) [��(�:�O�t X��_z�%;~+
����%�F����y��A__k�cqm#v�c�	C��!�8��}x��ܧ�����%��V����cʲ�y�/�����nGƀ@m&+��ے��7j`���QH~$"�_��UD2m��e(I����"����he/�JC�5ߙ|+��S��L%,Ĳ�	��v���H>H���|I6��|Q�Y�)DTd��ĭ}Y,#~���2�櫣�VXp���U��!%Q�L�\�pa�U�p�#*Ue���sx7���$�C�r8?M��)��X�<�J)]����������\��8ȻBվk� LM�%ߣk��h��Q�i='Q	�b���s����*Wo�R]í�j��܍q�(:�Q�	(���c}��1�*�|�&�A@����T4�i���l�����j>�o��L��|��b�����r��v���� �~}�>��yL��C��SiO"QOӛ����ţ��E`�:��_2�|���k"�+g>W4(-�A��1�%�pM�uן�X
��dC#�ϖ�&�S��0������{���5
���FSE\6pg��Y~ Vxï����Ȭ ��H!��{R�5���]G_����%%7ɯ
���S$�s����/�/ȟXw����P�x����6^R��p�#�g�<��p�fc�]�f3����4x8nW{+ X1�"	��Y-��2]��Pĩ��n�)*�f��@}��;Y"L:��kj0F(�%���Q*��}�Ñt>+L��dw��hB�.�xEH�h��e�D'�CRU$�p:�^I� ʑS�7������%C�@e�LطS3�f�Q-�ρ!��!��#C �o&�R�=������r��5k��^��?H�ȝ)�$0���o� �(���J1���N&��� �`.���H,�~����q
�K�S=��FW6F+�C`T�$t���	!`�0��@�\���$�,���:;D,&;�@,��!h���ޕb0<lO�7�s�����T����zx��{��C��z�I����%䤇1Ek�1��aw�SWm�|�S���Iv?�����
)����7Kα���و���=�
��k�#T����e(iR|_9��P�Ng�.��+:��g/-����u�;�'C���=�[����k�Ơ��S�S�'����[��K�CxB�G�TX�K���³̭�`:�V,���^��*d-Y�yD�s7����l@ �#�m4V���9�{铌�]����j�o����u7�I/��4�q�*5��b���r�k�i��L�����ܔ�WV�l�J��Ƚg�\\�'Hn��Ѫ8-�]�����5^��o������.x�*���0�zof��6�XoQ��U��f������6� [8J���9"v���lCe����A�97Ɲ�и�u���I<=��	�G��O��f��'���)�ٯb�R�SO3;���ެs��KE���oW���v��p�.�J\W��m���h�N�� 9X�71g�d@"��<\+�=(�2�}���~�|#ub+!�i��_t�������K�2�>.pu�C�L�*�w���"b�>�M=�0:��3��3��4HdU�!?x������X�G�oR�zҳ0���5Ĥ�P���#R�q��
9��������#i���l#]�� �NM���
ڦ?#j�>�	��'�= (��*�6����;�D��!�����:U�Q�ZGm���c؜JTm&h`��м1����y�69���&ȜV�a�ʨ�`@�V��{	}wD���6��.1�;W^Z���l���-�����"w p��d��4�3��P�߅e�x'���q��[�
<WAy�5x}�]oVf� �_$W�=^G�"�6C���������<O�| �\�8%������0�|�9 ����	�I��E���+�9(�
� `���i�XB�B��cb�[���HX����<�]�� J�zYr��6^��UX�ށ9�G��j�Ke)���eŊ0VA���&X�
R�I��,X�Ϭ&���iK��o���S��� $!�o�'�͠X~�͎m�����&=��P�2�ۙ̓�ݔ�t������ﭦ���{���a:����N�]�m�Գw��~�������{��i��6}����񛕎��	 ��1Rf��Sgyb*?"��]�k#6�Ɩ���m8��O�b��T�����Y�L��)���~�vu���Y�7��CByO����9420�Ϙ[��ߩ����ռG=���Ϲ��Ph��3Uz�'���̪���`(N����'��:����DJٝ�k0��ju�����RP
u�����Ԛ��|��7=zCJ�c���eOb=	�.����U��������ϡ|�7,�Ss��Ss���#�7���������kL�;B[���2՝�0V�m�\8x��\���J�E�l��i����$0HLCt,��#[�YvE�.�!f�J���]��H���m��D���ٌ�v��&���d6�P��>����Z3%(�2��ܢ���}@�q1@I	�QnW���A���6�4+����d���T[[ycJ2�z�-�W�V�� NU�jL�&Է���l���j+i�#��)Sa��_��m�N���]���7��=6-P0-�@<��a�z��3�݋�D�]t�S^?ye:�/�V�������Vt�d�ݥ�E{�����"�-�ηsqw��t�W����'��D���7�Ή��@u��*߅t�Q}]i:��~��MO�4���'�N�/Ǒ��f�X�[ �i	hmitDO��W6J������|�����<ӟ�����*��xoi�)J��{(��r���L�=�3ĭ��kF'��%d��,�=����vm�7�ꄲ�M�<c�wAS��M��������00�D
Df����o�B��K�¢��Q`�Fsr�m����7��ݞ�We�YAxn��@��{�}�EN\3�ァ�HN�W⚀���z9h�t�k�c÷��\\��<ɫ�O<^ρ[�,yJ�W��*ȫ�CH�M�Ǫ�I�4S�g���hd�?�ق0d�@���Vq�Pn� �%��mlÌL	;�o�����gA�D�2_�Pt�����9Ʋ�B�/�X�Tum���-���fE3����?�4����\T�_����Ŷq;�x����3.I5���.��\�{��".����s̓��-eC�+@E�_�WD�:W�i�c��,��T�W��b��!U�i*>0;�V�5ᖤD��q2��� �Xm�&����Ҥ�3�����ڰ��Ė"h欫P�RfU�)|5���x���`�൉�~�kMk�cx��K7[���̉�'�[���y��J �fٳE/gϧ[����5���m���{�Jͪ�&�{E�h4�	�����Bf��Gz?��[E�Yc3B<��5PY�+��%�'�\4V���0WK��U_,�i����۞��;���h��Vv�]�҉����[�u�W�Wb�A��o��]�qh9�}Sn��<cF��$bof�?�����%�
���~,��i���^�3�:s���v؜C���R���<o��XP�2=J���2=��b��O�#0`�|@�:�7���X�7�q?��Ǭ!�?��ږ����ӵ6��>��d��1D�f�RݪB�
�u�fbl��dD�N�_·}<�P��Δ����=����,�R  fO}#a��\���ҙ�)E0P�>f�#���x�|��R|p���8�R�B��YRZ!��z9��[<�|8��{�9]Lp%F�+k���r��h�nq%ڨմ/�)������8sڵl�p���xe��Y��R��n��h��R��S�[�������}rI�.����&��>Q�0�a9�&�ֈ�/'���)=X�Y5��+��;�J�o������)�Q]6�UƸ�6������=�;tQ�6d�aO���l�)�F�p�f��l���؜�CP��4��f_�J��|$��~q��LG9���>&f�C�����v�H]j��X�2bK�����f��E���x�M����3~�DH4�$�l_������x0�Q9�]Q^bB9cb�L=m�|D��v4���g����9wO�z��32��]�A{~�ҋ����t����+���'��AP{�9W���2�����~}Ƒ�)�&d彰�Б�@:'�c���b�32�>����I��+��H^��Q�9�论K�6^�	���tI4� ₒ&��P�|��.(����B�B���t�˩J��#����l��l����<�l$%�J�vfx��{��Ž���}�7�"ֶ�ろKކh�yWA��M�۟%��Ϫ��UYj�e��|R�$���NC�t�G�Q9���o��~]������X�"N��H��K�<F��;���`�"�����@}���2!"��7[aLec
��2��.�=2����VG�bɍ.Zk�	.�0� V-
����ⴰ��C����"���c%��y���X�>߬D9�=�rL#�%qEF�y����fF�����Uu*=�g�^�Xcɛ�9���5�@��;f�g�ؽ�������T �vc�,��|!m�`4 ��DJAf ��=V��`�u�8d>Sh�qԃP|�(��
��%V�ko��X}OZ�\Y�c�$VBߝ� T���ęl$��a��$FQ�p��<}ҕ�R�o��������g�\]��f n��s�1v�+V[jH��:eܶO5F�b\L-�rEj*�y�t�{#1�����Àu%>쪧�e2i�f�c���+i�[&a�f9#�G]����B����CЩ�BP�R��T�̱g�H�٫c�&I\����6t�����C��Ԁ�f�ú`�������c N�M���.�v����"��f�S���Q$��O����x��>y����g}\.�������@�]�-����2f�pzT�?����#Z��֖Ax�� ���D=��,�n���gUU���9����S���q�F��#M�7q�\�h�(���/p�`d��H(\4�j�&�9�� �U䕭��w�7(���a������?��F��R_-�4�YzJ�^g4�����~���@Ϝ��^��H���)��#B��4�)���d= ��3�3g����
�j�Oл��Ü�m�?�1�9F��/��@���Z�+��T�8����ط��^֬�t���ٖǇF���������u��^�����d�섲��s*,d�2�w䰲�FI�����a9���+ ��Ɋ_N3|�$>o�8}� @+�"j%q5@�;Zf�j<7���D+6I�,H�k
ӧ���@�g�ut~���e�!��t���).Z]�K�
��1"�W�����G�se;j�����t!׵s!�v��HÒ�PC�x;ʰ�ڋ;���?�|��ۀ&�iVF�M)Gz�J���03q�+a��N����x���A���1���j���f6�X�Z0�7ž�Ue�>��,���U�p�o9Ly����A���`��X�t��s��\�&��؎T��9z0�N#ݎ7�Y�73_�jm\�*�
$N�IL911�	kϫ���w�����-��ʶEM?;��<`D�JI�=bO�pKQ�mѽ�f-�3��"D�E�𫃂S�#6w'���21 }�+�kQ�<B�_ZYF�5{s����c�
���V��ROuS��H���!��j�!�3
{q7��'�EU��	ǩ�GF��Iu��Vebz���j�qr�e,�ܾ1����6�@`�d���=�n��Jr�qҭ��;�=�Yh���A^�0­}W�d��n+�B&�#!B��S@����b;ۮ��!����_�	��(��I��LǗ�Zm:Y��;r���eˏ /2N["�l�yͨ)���5[J �v����s�Q�3�G�y,��ki�,>~I��G����ځ�]��o�2fyܾ3���,��+�¡���8�i�%A�\�F۾�2O~�I�����F���<n�N��N���CB�����Z��Q�ҡ4���(��Z��G/�����cQ<�.6�hS;Kɼ����- �5��,H3׮?ɵV��/�g��%ϺA��v��#8��t�D� �`�rz�W�~[刎/��x�$*g'{s&���z�/�i@��A��i�k7�dHa�/�nE�H�4;~�0�Le)�F̷|���i>�ҼQ��Nx�u��C�����̽���=��HƯ�R�A6WhU����iݩ٩`����bˆ��m� �H�Vŋ��z_%�^�tt�Jz��;��Eԛ�j�Tq�8˔�K:ukў�+uV~�nA��S_b����gyC�~P�l���4�Z��h"с~*�����C�>��k�\���n�zO�E#�Ծ)��S�{�f�\����ߪ���ڶl�/��\��/��9�R��x.C��9��F)����%,�s����D<�%u��d�@Yf�Fk�|�E52���I��͖�`?e����l-�0@1YS�*=�<���B�5��A/*��}���Yr������U���q���7n�?�14��� �G�=m�^Q�R��	��Pύ,���;��Cq�];�FSK����S��T���5�-S��u`1h�S��+�C2��{�xQ���U,�D�[O����՝���¾�
��3F�`3Ӣ�����>J5`���|��I뱣�=�^%`��׿j?�v�NN�!n�|3�f�`�%2fA_/c`���Ҵo�	Y���2C$ڰ'���Ñ4���J\ܺ)��{$��m&X�����T�@� �W���S��k958�kR�����%�7��zO�s�*7��E�K�R�l}plLt��5��0\H+b�����0�/Y��vឳZ3a���zP��;��wO��l�m�p4�	��!/8&^i�!	�tdD��3�H�tԽ�.�d-�<�D��C��'o7q�\�DN���T���;��q
�b��]� �>џG_��EiDXE�能�%#B�
�lI�-�:����F���CԶr�{�j��ف�͋qB8[����}��K�Z��_h_م�b�}vLt�eZ��ͤ.��OM4{T�f�\&�:��Ot��vG���#k,�������&(8mr�7�E;��������A�No���8����*���b�r���=�-�#�V��"jm����^���?��QvW�n�J���0�C��t���x�?pY܅ɻ}��b��d��Xm�����ˆ��-�N�ڒ�7�)[���K��`M��7T��0�=�WժOF@�$e�A�0���rNo0��3��H�ƥ�g�(X��� 1��u�-�/����͕�Z�swh�e�wE���8Z��~��k"��oKM6DnU�������pB�Ɠ�x�S.�m��ӭ` ���� �̊�@C���k��6$�㊻Υ61��!6d���$&��I��������}�?�<��.T���a�[�#yѲ���ک,� X;�UXՄ����SH�O]�(`��i\e�5���ƊS2�� �fQ�#5b=^Ȟ�P���l�l!�
�>���-�h	���Z��V�Bw��A}����)�&�C�=,��T��J+4��j)��#��:B�0)й-�v�M \Ȅ���VR�"�RN^��G���d+%w@+���2}�o��nM14�������"i[U���^��U��5�?�l��RQ�8X�A�=�p���kmpo�C�I�,�gS�n�Tl���FN�O�,)V!]�"���g-JXs��"��I�]��%ԋI�����sU=�a��^i�6ճ�~����[_j�]�AE�?����v�/��qP�#}�(.�d���ovb%)?����T���h�v_���P���\���
t��;���k�R��.��d,8qnh��>�ϐ��f�ۖ�F�}�1��o�8y�L񚀢��jX1�6���Rc�b�[��U�rJ��Ze�j�sp(B>�r���u��4�� ���3�����P�3݆�׹Q���T��0�)�6�5�gئ��R��rR���a�mNS�����b�m�l������ʶ�K�Y�ށO�$dX{�>n6�z��JQe�%�{E��6_�O�=��#��p׃"�&rR`!Y������"Y�<$W}�((����.�`N}�z��v��W�CR�J
���HKMo'�/NL������ET>�~����f�f�`v�����V�����&RU��u��8���7\�%�\đ��
"�Pr���4�I!�n2V!�O{�)�*z8�4���JN^�h�S�6��u$�J����w�{���H��7(��j��"�3���8�s?!fk�z�^����x2����y��@OJ*�Lۮ������0��0���@�vZ��?F3�k6�4/[��� &���5���*�IUV�\[��-��{u�ғ�؛>�j��o�:�<4}h�u��(�O49`U�	�㽥k<�~����: ����ϻ�=���~�E�_}S� �
�����͚y��lm�������/��NK(L��������m�Y���o��.��y�,�jUZ�o[����W/Tf�/�n�r��;����@�NaŇe�õ7εCc�P~n�L�XN���w�\�ؑw��E�Vx�/W�p��͝	!Ů�;�4B���]v�>��P3�?'¸��+�!Q.�7g�X�3�����m�1��s���s)���������+W�3d������+�M�!�,�ޙ�4�p�_���$*$]�6|3x�9싡�]��)�!;"9=��R��:``��F��}>�� �1k��00�d1��Y�~c��Jnd>:��o�J�����h��C�h��v�@w�&��ɳ>�Eo�m6�Ala�,��%��>ե���E�0��]�*������NO����F���!o�(�ʊp	t��n�~���� �YO�N33��rB7�,X!�TN*q�ᓳ��� yK����W��.·x?��'pJ���%co��k�gA%��yP}zg~��AM�Ta{z��hN��S����j`�yDN{ZS�\-?�$��V���M^�x���>)(�Zw�]u݃����C���CJ�7_�ٝ�Ʒ���c�K�ٕ0���I�D�)4�GN�{��s�1��s��f��h�5�|�Sm��SOv=i�L];����g�6������>�dtE�xWя�{<�t6�����2���KFb�c!��p��r�{���?Ƹ��Q�4���~��Վ�',�N�^{Iogؘ�?��{[����F<��#��5Rx��aQ�x�Nl2��Tl��`Bk�E�)�Ϟ���ۼ:�נ�A�6w����hh�M��'�Y1�{�?Cȝf+��̭����������o�ʏ���OoKL��A��嵜͊D��d=��ݐ�.U�M�DA,�ڲ�������aT4v��}��AR@��.族�>g#��g��͗��!����c`@������Cm�9���Oh9,n0�~��JO��s��&�hF�6��no��x��i�317�I��Ca�]��gx�����kJl����Y��:�;�Ae�%�Џ��4@'��s6�{G������|'F�r+u:�	�(q�t2B.�\��,�$x�`a=$��F(sWי;.jnϪ�Mn띩��)� �i�f�Q��Bܷ�)�|�W]�י�"א���B�Xn2(e%~���6�e�eoksx��V^���p	*AJ!!8�)�_�>�l�� 8V�nu��a3-	��r�6�yA;m-�C+L��Ǳ��^I�ӫ���)���&�;��uݰf\(Z�E3��|��� ӗ�"��y�N��Ζy0���ijH?���[W�Qo셪����r��p�����ÛD���O��>:s��7��E��#%�_���?���%�q��f�f�4��*gh�	�>I�g;��� \��|`N'�����#/����������)E�ɴ��Eg߬��4a+0Þ��)М֒'[D�rܬ�R.�&M�Xл_�AV����2��p���=pq��.:d�ec��Dy�Ή4��o���𰕮�`�ګ�dl;���^�b#].��<������Y�3�fr"[N���&�d]��qp�3�{�D���Wzk���^r?*�����S�[�f�M���&A�ew����#��ӓ����#E�2�ɋ��Y�%��q;�W7[OK��m
�,����ϻ�O�k}�s����r�E��1�Н�O��O" 
�K�H��-�J>ø���,CÍ1k-�K3�PDY8�v�	��R�n�C� [������
�x2c�:EOۯIE�k�=U�B�թtq��/rQ����[���\�|u`�T��Pk�E��ɥ�+�ѱ%��H���;ꤾTn���  �����#��lx��>@/��� ����7�%�# W��=��o�>���.�?�hX=�B��D8�4�QN��``{z��a�`zi��b�[$��D��*�9�^p�a�;�nsN�?x���U���=���oȀl��ш7�����^���tO�ךp�+k�<��#�m�+�2��u�H �̈��g_ܪ).V'�(Ⳬ`������f�Z_��;�U���쒀Wv��3v}&@��Nb����롕��I]���Z-�ϴ9���z����>�u�PE�R�+?M�U�xf��BS���@� #w׬�s
*{q����J)A�R�M�g>;�>iZ��	�D��ENp̾�،�R$o_��s�PR��o����U'Uh��9	"r<�9�j�,B%'	^��&���3�J�~3��P;z�c͒�o>�h�JC�VéyQɆ�M3S:l5�%�rU|�`&HO�(~��$�r��]K?g?D���Z��{��MG���עN)�)I� 	�$�����4����7�v[��V�:��>)�x{�����A{į3 ~�%QԼ�/�w��!)�NЎ��3<�h ���8��7��lX�d��sl��k:*:иI���t;>H �A��X�4�2����*W�P3p^�B������V!���P�> �ˌ��M��J��$�m�<��Hf�iO�?�q�w.������ar�ޠ�����M�[��M�I8^@j�7��eGpDH:�}���	��� ���ޞid��1�h��{�b6r)��k��P�Sr��j&����.�ƙ���{g����x�Zl_ڑ�^��-�|p�t�C��Y���M��7޸ ^)�BTJjP�tS[� �v"��n�0���8e�څ�=6�3,��~`�d?Է\A)xߵnB���c/_�n�C�ä���;�g���9�O��Gy��U?|�8�.<S���xJ�&�p�Լ,�Q�М� � �J���H���p��Dp�#�It�Af9���r�-��w/�Ck�i��
��(�nv�l��)7܊��tV�lQyYr>j(�4��!���v��@��-:1��d�ކ�/҇��=��_ф��zδ�u=\!<v����uk4��3u���xl�)�ge���H�a|F-���zX�ȐF�a*s�[�uD3�|Tf�N�|x�sxԫd��jhKLwi{c�9���*�b��k1��ӣ,��Ώ�s��hQ���͢�ֳT4E�'q�w�v��4�y��ln�A�v�VmI��z�[�h٠5 �b�G���
t�j�4�s��V��{J�c�&�V�u6���
B���7��)�hI���v�������l��ŬLw��$��۴��쿷F^�#;F�9eF��|�6�FM���e
#���3���rh~�*��*^�����>ѥ��7�Cx7/y0�@�ś\���I�!�����ҵ�%����>�N��ߒ�f�"���\��"�K̬E�u������b2k@�I�k��m�b<8t�<�Z�Ur�����`��G}M+&�!`UtŗaE`KG�>ژ>�Md��9�&��f|�"��I��˄1Ŗ�S�\�[�����j'*�h��0p��]ӹ^o��<g��~E`H�yZ�ˍ��o���jXܣB!9&w�dU���ǫ��#����:Fѷ+N�
��qXء�ނ��wT��4`޺��q����DU��ߝ��FJc���C4Y*F.W��*��kd��P��h�<)�,LKK\j��?�e��
ʒ\����A�:�����)g���4�7sr�
��
�1�Czwm\�;�w�lQt�Yg�:�0sS�d�C�Q�&Jz��ʳ
/(�+1�d"���;`�C� t���5�NI6�a����@�Wb�L=7�7p�l��}QE��r>�IQÈ!CK�=�~�U������>?��3L{�7;@��&	� @�=谷�0������S:�f�d�9�S5�d�IgցɤdƠ����	>�r�ME#P�&�qGnv���6�7��#����/��e�p+���'m^!�i�J-�m�_�Cǘ�9�U������yfQYr�W@6@d2�%��m����`�>����h��(����g���òRd�����!���S��W�q(�F~�6��bd�9�Y�F��;��4L�=����6l��<eD�>E2���pv�] �,�����=eP��Er^��e�9���g��b�x�4#���/I�D����mt����<�<V���;����f'�!���w�[Ap�3G�Qs��cX�w�?�>�C���������S]olo��H��� �R.��>��<1fG>g��
[� ����WN���\����G��[�5��.<03&�s���^;�Li9J���CO�K9H��>x�����B�d� ��@-}ʥ9�<����Sp���iR�׵�罸�(Ixks��b�%+�X��c\r���{�HZ�t��p�&� V�����:F
U;`#P��vS��3�����ֽ���K�L��i��D�3�,ܫrx��m}��%�_�b���{��S+�@�הT�c�*�/q�셕}�`���A����8��8Pwg�	�<m�Gs���m�Gt�w�Im�N `%�.���+�+���l���L��-�c�=�X|RH5rJ$?A�~]M�y9!�����dEJH>�FL��:��O�[l�;�b���ҭ�rOKU1�ܳH�K�s+���y-�!�q2R���Ϝ��Zi�%��=��x@` F�'�F�����vE�[8yˏKfoVaV	|�;�!�wfI��%�l�Ó�tq��횞�?���"8�a��J��\��0�T���&rehx��v�e�M=8�S���.�-���	�e�_�0Ay���P_A���x�y�~M��2��j����{e#_�ǋF�]�������ʱ�K>6{�+�����A�!��w6r�ǘIZ�<�j�-���p'�M�������{P�|xڬS�(b޸�2�B��L���	7�hЃ8�|	���`�LMP��/��tO�vO�%��@3PK���JAʷ�Uhc&0QL�A��"eX�����N�i{Cf�r�x�>.n ���(I--���W�/���"�/-��zyAo���t�/�K<F Ŵ�<��9,�߽���.WvTyF'�%���Z-몺n�C��V�&��/�y<�smM��wef��&ӣX���)x3�GQ�E��.OS��?��$V]A�4����wR����[8�������M�]v��ɮ#�� ��#���n����I֊�:�t�:�uw�^��>Ò��a4�� �_�fW�28xFH������m:V����@T������!�8[RL�Q-1x��:^f��'>����&�mG]��E�m�l�<AxK/+���C�L�ԄgRxmeC1�+�\�T�yO�1
�Q-�s����5uo�`k�Uo^P-��į-lec�t�@0v�#&��F#����9�H�.U�z��d�=��[Љ����!�'84$���ྥG�O��b�rY�p?a����q?qp�U6,��=Gagc�N+�"����+�j��J9p���5z�f@�.��7<��It�vzM��3�ǡ��YH0Iɪ���Þ�{��fw0� gr�g4�stȢn��S�5!��IɲJk�J���r1�"�E<p��d���
X�l*{Ђ���4��͟jUis(Hj���>T�� \)σ�!ө��f@ȧ�b[kvE�4()�5��4;�+�I��Y�p��K֜)���V�&����e�X�3=��!+�,�ǧ�l��E���b�þ0Z�X�Mj�޽��nW��P����"�J�-9*II�3#�#+HR�{�G���I�6M��MK[���֕#�w���"�@Q��@��qƈ���ޡ ζ�ÿ"q��(���_�x�c�r�I�*�Uʛ��P2��u�@����QD�ڳbZ����l�� �SV�NÌ��׌(%��bb��є�m��ZKC��X�r���'�����H�y��JT��41��dg�d�V%�u���X��%��f���R�p&Z-$}xMϛ�_���[*�5� 7#�*�����?�?j8��?|�:U�@�ZgosC��߇�)�����)N�J��A����8(
���	æC�^������O��3�ݵW��qM�0U9瀼鄜�fx2�J.��r2�������,�g�{?�|Mzu.�f!P��O�b ���&�O��].����	5�b*^�F��_�@e���*����R8�z6̕h�D_�]��*��Ȕ�nW��_���-L5����0��z�4���Kd���bV�����_#r;Xbc����M|�[����~���T����;5����!����2-#�%�N\�{ͷ[9������	q�|*�F�֕%M9�51Z0���/ds�=v���a���_�!�7S׈�B�u���� 24�R
p���,�ŭ�VR`Xfhm��G)Zz�K����=^R5�lW�3�5'�>;�i�*��3��"Z�퓐�o}F��&]��Q�K�-�c�r����`�Y)T}�V�Xy�sX� f��{qj����L>ŅZj�W�Ŭ��4�V�K*q�cPӂ	�w&�=�U���&�f�2	n,���&��R�
�u����oM����bX,�o��wń1��edwWM��%��#������+jo��K
�ËW�3�i�A*^(]`�va��ϳ�D��GtG���ҏw�]�"����]Қ�_��U�Ϭ3ы*����dZlY1xUKOhagp�MI��\�_M��w�B�5%��!�X\7D�d$M��걛)]S>�dgf��7Wl�Vb�
�}|�{���h;jm�����X���+�cpq�G}�;i�U�6��Of4������\!!9l�0~���.2�`�Q�zC�fg�4uT��S����V�Su��\y����.������H|���������)'�f �����bߛ�zȚ��Sc8�Zt����Րh][b�$xĳ|+������^����0�r��RB	�v��X����Hx��N�p]j���E�o(d��酱��沙��u���aE�4+�nq�}	����Y˧����Hp��L�薢Y��{�P��FeA�7	 ��s��,W���Z�Z��,�!> bwl�Z��������FBh]s��aQ�Wk.��W�P��w���g�L|�����[��E��*�=�5m8�mΣ#�c�P��<7�,��K���Y4]`���M��	�R��'�1����/�7�^�M.{7�9x������9ƞ��vg����
��w��{8~>?<Vǎ����$"d��b�Y�����:�������Ϡ�~6%L�F����<�~A�~�%�'Đ��������5���t۲!�I��By�+N�s��ځ�y��Ci��*PN������~���PJ��ֶ�[TD�Fam���vT1!�0�D�/��ۧ8�>xjd�ރ�'�3K-�����?R#e�+��:Ls�;`2u�f���Iq���v���V�~Hŝ��ٺ�4�y�0�����3�ZD��ՉQ)��'�����fY�W(K�#�^wv�J������'���*�
'g���v��
D6)3Kދ?F�M�����v-;1�$2}#�cҽoyJ�O��ٝ��a��]��Z�_خ(�hĨӑe�c�����k.�|�]��,vɊD֐�v��"����Hvs���'啹~�T��]����un��K*�#�T�P7g~|Z�·D镡��h�qK��ݙU�ͻ�5�p��Jс��aj�.k�;�����	ܔ�A��<��w�UPN����6%B_Ag�EX�����[�͍���tE���>�K����K;�}�*�QL)1�)�7&U6i��~���O�*��X�w�[�c�1�C�	j7G��=��\,v�����H����n¼a��e7�vp.�������%дV1�+��n|3RNQ̳hdw�:Ѣ/�th�g�;���8J��|��6�פ�c��>\03�<����\R�\ږ�G�����*���8~�#JNJ���v��m��q3���Vt����I]�~}���(�o����4���'���`r0*���F�����Ϸ7�KٚpNܰ��QADk�5��+E��Tf� ���W��\��U�"�`q��%���߿����97B�2[�n7�*^�idR֚Eo��5<�$��V���Xk��(�(��A 3E3�(ѣ�.�k�O�Rk\{�@Q:�������s��s��V�{�`��ߦ�F��9mݱ�����7�\�B�����3ht�mh��P
�u�؇�� u��oĩ���s�(�6�?{�"���)yk�~��$����(��ЏK�"G9��U4s���[67���8d�ъ��_���vS��#�Ew��O9�ȵ2���kz��a*e(�h��30�A�H�/y�;e<#� XA{�t
z��P�u�x����'BR�b
"��ǺOP��.��4Z�Z��*n�Y/�y9%�����-�If�˸�W���W�tP�@�lA��Q<��0��B�2��4����6~�b�����H��22����{c��u�|��=�vuh�����DƗQy�t�F��?���)�z9x�ȩa���4�w�P�����5� �����N��y:��}��	+��O�+g!{���TI*;x�~���J�ݢkٔ�
V?~Z�Ѥ��wSH�U!�}/[w����� �U!̥�ׄ��1{�'����SfE��f�B9w����kM�M\ғu�$��,�!�Y^2�*�aC+�����E�Sx'8�P�>���u��G����C�SaJ��w���VOB�IA6�}�_���Cv@2�3��u�%�a<������@e[s�x�M�K u��d��.���%z��
��)���(j�M��-0��C#r\�lS�V�x;NQ]�@�}�wa��S
��C���m�z����)8�.�0�^��mw��De�qK?�s��i`J�3������/���X���!�߫�lS�l��A���
4�
��H��	�����ثt�l�㰕�	!Z3a��=y�j��a�m�Y:�CL�|���c<����:��Z��rC��|�gu��ɾ}i2�=
-�w�O�)�`�ɕ�X29�~��h�"���?n7�p��a�رM��oy��<]����;(�!H}�yK���u
���	^�0�����7S���y�BB�� ה��Rb�l�O`MT�Հ/-���׉�ں7y��.�K����N���
���6a���_$��b !ĥF����O@�ùߝ�2q�)���|U��{��y�lۗE�E;�V�+�.�)�Qv��'4Y�N�{o��u?	��́�6��?�P�a��,�gİ���-�����,���Aƺ]���ӫ*�Ж]��,&f0<M�	�ܨ��]qY*�_�4l4�������8$�{o'L^Yh8'x���5��;1��Ǥk͊����Qڰ!���@�$"�b~��@�D�$c����{C\Xtw�w�H��ĉ_�M�?��5n�I�6���.Ţ���`�B���,ļ�2�߈<x"SHHK� ��'�_���,߼��6���6G�A� �Za#Wt�ڋ�7����A�k��5^��c��o��s�<`�>�QY�C$���CNZ�R�|�%Q����R�"�gfִ�,L����Q�F�X�Z��3T��(�"XV؍�<J�N�V[�����)4+ �Ts��;�;�L��[W0Nf����]��>]�o�ޭٗ����{�u�A�m`�h�,*�������P��y�I�C �~�wntx��i������g��ʮ�dó,�{p��>3��=t	������X:Z�|�z����L�/1�ݶ��U�I�Vx�Kg;	#Ez�y�H�A�c�.����Ӵ�O.E��� ��9�xכ����a�=���s$�o���6���U��c�H���:��H��-�F�>��	��<6���.���ߦy�[=�>�5����&-�Թ�\R�׌���]f06�\�IT+x�j��m7.�����D���ܗ���?���}�:��Q���= ����ߤ�?�s&L+P�nX^����ioc_7��\���8w�2�$^��o�(��������Ts�6�t¢��J]��ܕ9�F,͐�1��1��v�֙޲;����`�"����+O>[���j/sudB�'lDn�Ď��T��Uq�ih�>K�xi��������@��c���Nl�+-��;�2?��e��'a�$h�A7�7��a��k�*�ߣ��&E})��v�2a�γgK��%1D��0F��tM�bD�����	�2�.�\��������.@c�l�4vʹ��FM��}	�g��)n�;�����!C6�V,V!Z\�6�����S��hOY�E�c����+sD����6X���$�sҰ�;NY ��@���^֦���3qg4P��qdaa����@�+�3C�b�fʨ��ݷ�+>��Kg[j1��c�m�"DXSg��%�-3<���os���3��"�DԾkCt��-������{�&���eU��#sMȡ�T%�Ӭ��g�pC�h�	�@��4���{�=B`�5Bt��;�D*.r������^�R�g4�;ߞ����G�%��,%�.�*�H�M 8�Hv�Q\q�����C!$�O��.4�_$���؜e_�����y��o���my�K�a�E�R� �]?q��{����q�"|��q��� �.s��7��벡��� �{�	Vq�N�`� k&��4�9ͥ%��q�h�5�F+?ʣl�30!ǉ�:$��Q�n&��I]�c�c	�{؟��j<�����X��.*8e�³Z
�ӏvAN�=e�*vE|a{{}�� ��Ln��*팈�\�jH����!7Hf�
���܄�h��5������
 �c�!��ޚ�����S�F1+1-����&�3�e׽gKqs����6&DX��?=T�Ǿ^��^�k��v+����D���\�~�Jc��fU7�1z�#$;9�D뛣�׻.���e��
���+;AK �כ�C�w�C�����	�Wa�$���Վ�����>x��*��q�C+���#����@uই�{� ��fH+���7�r^�L��S��Vѓ2�͚	y�����
���Ys'0?��?����)�U�&&�r�A�����j��N���v���*|gHx 0p�����I�
)O����n��+�h����?�Iz�����T��g�p�d�����=cm_��LY��<����P�?̟����^���4�ZGݔ��)�h����O��}��������=_d-��m��E8�lR.�Dm��ӎ�K�ǧ�;J�N$4T���yC��%��|&��n�-��m%�+�G��-�Y�g[(�f>|ކ�Y��Z�R�b�MY!���a 񋚝	/>�0z#�:=��(f$ǝ�Ŭ?=��!y4&zx�� �f>e{�k�������߭b��c��z�K�	�SѥZ���ύ��}��S������B�tX!q{IgP�� ��B��R���$�Z#��ʆl�<�n�M To=��*=nh�������u�z�{Ǥ����R6amOU
���M���],�)��2m+�m��_�-�X���2=W�|��G�Y�\���������-��q8r�q�e5J��`7��1ꡛ��_H�b<k�O�ܾ�����. IU�&�3�8���5�A8�C�����'�o~&����MX�glͶ��4��^�ϝ��1C}J�ۇ�W�_{;}St䤿3��(c|oF�z��"&�[b��<�s[��Y{�=]�t�>����.�&k�>2�R�`¡Vb�F�����]%�ڡs��^�v���./�;4mS�V�t�&���Y+Z��*��~����%� ��U��	�l}�+{	�����sE�P6�+Ӎ�T�l%6�b����J�7�&"���'�+8F�7ci�o�n�=䑃+����A��$�F����L��	��V�"�R�%�sI��}�:�nG�r�E�\?���)�=g.�{�a�k<��ww�2���x�b�xmD�U���^���4j�'e���@`�,餧Ae�y6������ـ$�mu�q+B�$X%����9�:��lE�pj#;��>e�"��345
Z8N�.{�y���	�:�t�����#��>�T�+A�D�s��[��=��#��,����?k�����H<܆�9GڑY�}ñ<���o_+���-X;З�h�S�J5s��V���b�3h��syB��u��$v���p0�d�m$��ͳӝx�g ����_�B�<��Ǘ�gb�`W��$��hK�Nm�&3jr��
D 5��N�:*ۛ����p����"�qIٳbv�H����db�R�#��+=�������4H
����k>{_��{�?�~�'�=�����d�D��`H��껆i�'��y)�=*}�V&�L�"M�x���k��c��\����ɒ�b�Ͷo�Co~������:�:�W��ZӤ�Y�s2�/������g�}�ᔟV�&�Vz�['P��p�����X��h�Pw.���m��v��2��c]���'��Z#�Z��ån�Q� ��+�W���갻�͡L^X�'���i�m�C$\����J�C���%ItҬRl��;*N�X��h��G-�('39�oN�I�O'��Pf��Ǚ�Ŀ���Β�O� *z��>f�ʐ��̞�wd�k�_��:S�,�y=�Tif$n�s�`��˖6(����/��|V��h~��r-LJ��rFF=����`��۸P��qٴ'x��)Ɓr���e�(^�	��tP;�j��k�cGk��-ԯ�>���oB5KZ�hU8F-�WMy �y�ʳuz=H8�
κ�?� BPX���i���5����9�R���)F�0��!׸����zy�]q�;�KG��j�F�+׼̜���x�.Ґ�,��Z���p��OOTX@VN���x�j��i�]x8i']�
�V`2��8}��a��ED=�����}��H�b��y��0;����t��OK����훮9CR�
+[��A�*��/Y�5�SB�%��'3>Q�Rg}c �3˼j����.ZG�l���b����݄q�ɩ��ӝ`̘ilV�U�����G�F�{;b��ʴX�,��Gz��c����&>;)I�408�Us!��E�}>.M�+dp�]̅O���n5�RV��������_ՑV%�O�ĝ��%p����6T�{�2`�=���[b5�6������k�N��h����yz���pzF��Efb��i�ܓ�6����i�S&�n������U��{����%����,�Ph&��+N/ z�,�^��Z���(���Κ7&*;�c���cZ"��Y�g�x�Xv�
 z���R��{N�C,p�>����gw�2�u�o+m�P6QA�a����0mrN�m��

�\vI��bKt��x�A�_n�l%=
b}�r��c�w9�bIC� ����F�&L׺��`B�\��Du®�@
���V�0�s�h�#���L�t.���I�5�ه�ǉ�ƴK�cFP9]��o��=I;�k���I��ݑ�Y�)wm���0������X���ksb���~-9�p��MeH�^�	���$��^�+-�eF��A��B����� R�}P��Q\R}�9���}�ȕtR�i��I6[[PÕv 2���;���ޒ��y��kÎ� ��^Tz$X���������Vq<�E��j�/]m�7��C0Q��oi�Z.h��ۉū�)��&�}60�ݻ&nn�"V<����?��cR�|�K��yF��ߟ!�R,�t�{a���W&Uٻ������H�}V`*`�D�h���Gv8Pp�i`�t����>����T+�d��t��|��Q؊���a`-���11�Bb �}�;�%�ʯ�����b������2`ʡ��z�/�`�x)m���K�N��U���8�23���H,�a�
l�c�&ʄ_����oЁ{I$��ztx�>��ߖ��x��>3�|B���+Um��f����$&VD�R�&�h�D�����pd�H�^24#o�©���/j���߲�H���%��z��WL9Ş�뚋y�E��b���ύ�k�7��!�fB���&���Y}�Dz�lf���z�G���k����bi�L�I�3f�s	yq�o"{�<��n�&��1�>�M�Vo�P$�n�\}ϜH�����u��L1�J���2�ek���Q��7	�ۢ
��{�v���&+A��	p\:5/0���@�;j-���!��J��*nڒ"�¹`�����=�q����|R����٭D�%���~Ъ�@}�F������闋��e�a$_����ӳr������K��ͷ70��ܖ`��;\P+��A�w��^&4>�*��u�A��4 �8�+:���ʋEB���D���Ƅݧ[�KߜB~���
���KJ��\&�,�g'������w�kw�������͏,�����M�G�����c��F���{qEx}���iQ#������0�;����܏u�Y]�HQ��u��b�kJ&$T�C�~Pτ�S\@C�i1t[H) ~�����	F�_�&�GHIyo��%�z�i?�.�{��x�ƣl���^���nHxOE�e�S^�J[t���?��aQBu��,צ�ڰP��B�(���e-�Z��G���1]qc)d�O��<�3dx*�2 @��w܇����Yf�f��ZqCk��tcܯl��~*�$�	�۝��h �Mά����'^�(����$>:*���[�(�HWLQ]�$az���$��2b�Ψ��1s����q��Q������S����U}meC�i�M��eeF��ģ�������*���Y�;+�S�K��՞'U�SiwH*|�u�}�gɕ`1�@Z9(xP�佊�~��X�`�(���܄��ܵ��.��8�{�J��1P@��C�"��J��d~���Y$�q���3:����{����{}�Tj�ѿ
3A����e~1�K����<ז\߯8hF�Ms6}o:��P����&M����9��2��đ�u[�Y��w#�&E;�g	/g����5�/$ړ��a#O֦JQ� �>��hzg/nR���Fy���R�
Q�3��m\�{�ܞ��(Y����7�h%p*YC�w�E�G�ԣ��aZ�]�It����A��l�5J���c�.�ԕ���dHۘ�W�+�ä�v n�*$L��E>��d���.=P���U�Dr�SȖ��WZ���g�a���Y���S��%�W+-m?�+9��/X�n;q�~2="�aI���fe
)��ax&r�噲���+���>����ԤZ�-[���?~E���1>f��PCݖ�&�ymi�[u>�`�'�
��3�M�#U	_�)��?�E��a��ɘ��`��@��ook9�]�i���'t7�ó��x@Wa�|x�qZ�Z0:��% q���E<	��'�P�iL���5�2Q�<u��㰼�5�X��{`�B�O�1�����C�RD�JI���F�zG;����3��CS��=�C��s��qcriR���0��(�}�u��Փ2%͓�6�����%(�5�'%���"��f�O����|A���J��Cj�?�=[��M���
�i����=��S;߱ q�X�w-PM(����u� $"�z�,:UD����j�@q��@Vcxjǹ�ƚaBqT/���Z���erڔ���� �����w�e�A!!��.��W�LH���n)���INB%_ ��h�~H�4��{ފ�ʴDL�G��Q�8��z9y��fTk�ș���x��P��/��>�p�7s?��^dx(��ʮ�Z�f��s�R-�@��8g�~h�y'k��^��q^�p�O�Է��e.w#����g�i������t_`L�$���9$.������;uQ�iFX��c ��
!�<��_�yB&TǝZ[��n�4�UNU���񦼆�<|��J׊|nE�s�p*f΀g��b�����nL���Å	�팿"���3��/���E�&mc��`ٝ�t��'�A�8)0�[��I<��Xi-��/2�w�ؒ\�a�L���(�B�o,E��z�������*-L�6��~���5�a�۝"�2&�R�AU�hă�>�or���0{Տ�P�oU�X�d���Ih��,4�}&I��缻���QT�iL�N�3�O:��3�R`T4e�v�p9��,��������*�` N�m�*��� ����8fz)z�#Xn���RT��9GM�u� Z®4|'0Jw�<�x�H�|��y.)�'��j+��V}�9��˳�������oޗ����-�F ����5�roe(2���d#à�B���u#��s]�ipx�t�?�u�ͤkH�cT�o�ld�c���3|�6�[F�]Id�l����X��OlI7��8��>Y��^)�}�K�}��\d�hj��E6�mWdD�\<�=�ٺ��}2{�W� ��u�Νd��2��X���7�k*�c�FpZ[&!k�Qn��+oM��-�S�.v�ӢM.a�!��\w���xX��v�Z�n�5o��
���g��l�7\����ϝ��פ��o܍����oD���"�-��P^q^��A�D/KU�ٶa�|�l�P��4�֖	�͡���en��G�'o�]{w��ܨ@'f��m�`���������[sHg�^>��g��1�(�~�jbWbe��Z��Q��.��^�P��d<�U���oC����i&"�����z��S>��&�[��!f����ZaB�Do��>���$A��"����=*���D�4k�j����u��:Q"H��R )ǐ�M۰-���g�8��&\#9Wo0eM�\v�q�p�E��,Z�0h,h�z�:� �>�A�pS�t
/m��A��˙XN�H���#�U�J�g��$��n��jM��Y` [�4��SiU?bַ�j�y��V�{�"z����v����l�N{_Y�BJ�h��-���Y6t�����D#Q����j@�7[!tHp��c�'S��G\|�g% ���Ro[y�	�H?���Njm81��Ih��/h�r6�i�3a�}T�:aY#��&�zk����WV7P����;�S$d�:���u��(e� �����=,�p]�2�C?� +>	K*_|��1���|ݷ�6 nEo��ҭ)uȵ��=!!��X�=@�����_����\z��oE5e@r�|�*�&��2�Pi�E4{`?k�����,�>�k@�$�l��6Nw���K�%ە�k+�-��yo3{G�H 2%�y��ڱ(M����9���dc�D�=����E[,��EȔj�����rxn�$�=�Rzl�Љ yu|�
�Ƹr2�8>��q)qr%�R�_�=�3%7s����1PD�+D�̘p%�M*B�W`��l���I+@�oʎ��q�	G9$�$j~���9�(�A-���J��/�� i�`�ܻxM$�Z�[7{�{7��B^h;���YJ|�<�FW3x��;ߤ�6���J�'yZ*�T��|�:8�Y���dVz
!���u��Q��_s@Ϡ�����y)F,q����X���_	���:E��:�%G*�h��
���'rM*]:A��@�p:r���A�(�.���������4[�닕�8�T2U�P���C���B��S��M��A�4Y�xy���p�����<������-�7���"
8����0W��*�mB�	>N*�,̮l�V��(�f�ɷ.˥C0[2okh�Oz������4$2��.�Ə�B0�	t�w�ʜ���Cs���%%���pUj��5Xt����_����'�6dR��m�C���#a~��_^�5mN��Q�>���ֈ�AL�uM���'B~6�+h:3��r���3�&��(��0�� �b�?_w���A[�[�� �,�<��Tj���>��[�����0!K�凛�-`��w����5�;L���$��xXU+�r�&Q�s���E�@x``������ߛ;R�%��3>TL,4�)�E5��4��"�;�W��斞��7_g�%�j���1��>�iǏg�����0����|�qÉ�]��(l8�}\Bql� ���(kF4�8������ |��G1d�_�&X� 6��n��fT&K�j����x�pl��=t$��(&��|lm7G^@=�X[��k�����ލ�AZ��� �3�5*6.��b��Y���7'�!��:ej?�U�i�����'e1����2����+s���@�D���O��;���r{����1����KġG	N�QrbH}*ӥR7��1��鏄��$[��t�,чb�7LBr���SD�
��$4p(:��~I\�	�ӈ��_���������cQ��*<�+�ֽ��Z��囝S��偁����'58XX7a�<:�R���!��Y1��^��7�*�F�rER�4Va:��ٲ�)�-�Qu�7�2k�ǆ�`����-ޣ�s���0���n\7��ߢ�Zp��FK�߲\���%�/3���7�dI�B��tRT���W��#�g��;�<�y%z��Okj܁ܬT�!ZR$��zy2�Oj��~���KRCLH��Ƙ@Ce~	Sj�g8�l���b5�08��Yн�<a��\|��F�E�S�q{y[�!p���tG�2lp��i�v"5"v0������E�8ԫ|�
��NQ�!EK$��HbcH��!:�y(��m8��3'�B��]	����#1	�ڿ.&��-�k�\kG��Q����='�1��O�p��Y3+2���о��k��T�"Ϳ��ycX��|�t���pvy�Xy��1*DVQ���`�R'��7����J�c��2��8堪~"Fj����P�w�k,2�����.��H��"YNs�����Գ����^�}Sr��n������t�>�2:_;�ּ�n�,K	n��7�e��Nu+D�;��8y�4X1�&��U�6�Q�R�+Lb���h�����Z�s��T��{"�-1�#8-�yY5x�:�w�??���,�Vd����1޲>8̦D��r�+3j�/gh�\������֐FsFj�»��\;�@�̧<��SY4yQ>�b �aK�*�����&R�%���U1PS4m�Ϣ����TS���Ԗ�Pn�#�U�V�?�`�֔��@���$�U���]����R�f�e�y���a��N
���Cz\�e5h�b����&�f=OL��V�(� =g� �\x������Z0Љ Z����nVU�F�~�Wq8�ӛp��hz�3���;��ZiG��dB៭��/���k+V���(or����'M3��d4o*������!�2'����u�D#�;�,#�x�_���!��&s��������>�R(����-%�FWT�����:FX�����'�1ͥ�S"�9.��"e�g�wwp#Я =1Z|�(��[�Yêg��6���M��b�ݛ���~v7��Zc�gڲU�M��.���{0�f��B�YҍF�yB㹭��3���w��$x#1��|��d��Ƶ�?��x��>�ݯ�o eV~�.��-�gQ�S:6k/.&��s��7�4�NF�%\*�k�}�	���w]`�6��=�F�GC��iO��`7�L�� `���k��<�Q�Xȍ�%�Jas�GX�B)x��@������ND�"�#b5��D��)r#�#\k�����LB֯}{I�9�Dz�~�S�����r�.�:��S�G����X֐��T;_�D�FV8�8�4�>�S�W*H�P��P��O�Z8�9�Eg�k�)�]���?��#�����=��z��:�X:i�~
~H��}ը�3�Α�Hk��$%�BwVm�.��\�`��h�&��v/4�X4�Fnh���r��63<GWodĒRk5?d�X�./CNOnW,n���B�F?�s�{퍔�{oU4��~@h�HL��ן�`�u��������l�_�{�v��ⰷSC��BE�*��N�˔�)���p��9���c��P�(��g�$�^�����C��$�����7�H�g�l� �LĲ���y����/��BIn�.�{:ߔ ��jZ�a@K^7��~��z�sb-0=�2�8d�z�5�4�xsS��7�7.ZLd�nq�ؐ��	Y#�M%5���]n.��=��S'�.k����̹�s��)����dj㌮mMEZ�tv�r�UlKw\b�ߞ�� 4�{{�i̼ť���e���Z�cp�^���H�,֞����<��̩U5|L����<�bM��qI@z'�+r<�I3���?���s�Q�U�]!���)OX��_s��<wD�Kά	�po|��\<���S�R2L7�de\�.ʫ

��O7"��èI�����UoW��ߙ���*����ٺ�f���ڡ�)w�=h-�CΓ��t�#������I���`�zp��q��[�2K�Ήrʌ��������֖!&�#�[�z��㛉�����#Y�B����W��|Z�MSD�"�L2fu��5w�eҘ7E����]�;-�}�k����d��fÉ
k��,�u�<��'�Nv',��Sȝ�B�x执D?�Щ�a��t��!BԌ�A��~Cx��5�l#�f�َ1$�>{*}p�\X��%i:����ܝ��ɘ-)�0iyQ <Ƌ:c����e������u�=���0�>��兹u.�� �����lo�r�����֐�Tn�O1�����ց�bG���ȋ(g���;*N�����+ �~�?'ד�����P�}�O.=�d�����oDE�L��$�߳ގ�UW����0�8�zd����3؝�硢W=�i�N0�x�1�����K����p%�0���塱�R<H�B;�]��c5���jKpx�t���� ��Cwp�C96W&P��]b�LVn�o�������E{uZ�v�e�:����[��jrm)1�e$��)u�&�y�!���N�{��[��Q��M��]��P�1;�؂�+=����Z��b&�eU`^=�v�������Z�c�~7&**�>�4��q6F�����4��&�:��l��X�V�Xp���K�/��Yd�xR��W�\��ϴ�����_*��T}�E ����^�(ұ_Q�z��!�_��x��g~�����І���P�U��a3��b��.�m�k&ca��/�$�FF¦�U��S[ěi� �V��2]&@����G�x�\&���H���x)��}Cf@�y(W	�iQ��WW�UV��@��ݳ����с�3�VpʯO�a�X+�{��&��+�D|�7u�~�d�UV�+�L��ʒ��uDI�P3@Y ya����|
E{� �< ?��ɣڻ��d�H������-���*�����x���{�;�!�k�iˡ��+^���V�����#2� �Bظ�>s�=`������Jj��af\"5������GK }kY�V˪��;B_?&���$�q��Y�Ԯ$�L(������4�
���Z��fo���SPީty����
]�l���>Y�eRnBc��bFzN���X&]`�S�0��ŀAE�G�{�Q|j�1wݙ\4��e/�IT�r���=�b
��A�S���*m��{[��+���+Ө�����ֲ�XI�fI�j�.�W�(�~���,���&�@	)��W��vBҳ�A������k��[�S.+�o�o����E����t��ϑ�H�ǃ��vG��a��Ж�|���}�ֶ�$�.��^ˉQN��
M�� u�g	�h\�(�\#K��^�Zm����62A���=���7t7�Mcngs�'�I
��PpS>���t�x��E�������Z���R�&�'�Ac oS���j�q�!�����l:I0�!T���d\%��Ph
����' `��`	���]}��T�F�,�[)��)�Rǿd�{:����hĕC�,��9wȄl����5!�=�q��'�Q֥���y��<�!��ѕ	��^ �u�U��E!�Е�$�y\�n���1�3~���B`9�Pډn�n
ODx��@���ԃyW35[������m��1����:L)A@G[��������^����$��.8�k�/2=�i�ID	Y��R�8��h��7���Z��P�˥:�4��7F��(�P;^�2	�o8�^["�đ�N�x����M�"c�Akݙ�p<j.�D1��@��3o)vQc�#�%o��3�ŉR6��Q�=��d˴�rӕu鞑��ؾ }�9��4� ��)~!���DG,st��A'���ӈ�@��`���β$J�d��P�V}<ʬ5�E���w�%���a9�s+�$j��h�/;o�hc���Ant���#f��ә���WFH�6W�Ƣ]����p�]xqd!���j�0�`������g���x�k1.�v�0���;����a�ŗl~#��F-�-)o�.P�Y��Y煩/�4>�&:�La���-��f8�G�{��KϏ߬,���6�I~5$��ŨDJ� ��y�����z`��k��r$�Mu70�QX�R%'YZLBep��8Ʀ@���ra�����d2���+����k7�-RΑ �jS=����Pѿ�.��h��SKŪ%�a�i��S�|��~�h���	��5j�� 09k"�������p����c���y����(�fɟ����$+h�*w��1fڅ�� {���6���h��pٶ�?�����b64D��),��V���"kf��2! ):��Թ�a�g;�2���@.��#�C��җY4���SD�BbCԷ�����-\�7�o�����Q$S�=<� �1�
z����k?{�c�J��C#���5_e�4!To2{�^��~��B�0���v�}T���!T��He� �>(�Gܽ�X
���v�TΩ�n��rB�bD��Ƭ�Cv6�cM썀��^b�%?�t�v;���T@o���Ei�*ŴJ�}ō�ʆ��H8��6��n���?Sɭa��u��.a�M&ڶ�l����.�H̠	���C���"�q�t��)>���o��r[��_��Jj��Z�:���7i�߭�-��Őֹ��%G�M�P*��*,Α	6ܲc��O8��+/d
�Ҥ����"l����8/@��8|������/��#�m�� ��6�`��",F��r��t���H[AV��� NcAP�ɕ{�+�ߎTh�ІZ���D��/��ع��W�e��k��*(���,���f!�J�N`+�v[h����oV0_��B���*�)���$��\�A����&���U2C�K�*�n�js��*a.��Э;_�9������l��ba�ź���2�o�в�r��>F����'����1褥/g*/*��$��1�a��b&n�H�J%��)w�?��z�����.�X���l�7�I$l}�|�az7����Yx�\��:��!�Fz���M����w��a,�$iF�S�=�I����S8ҭ��!�JS�2�J��xr�z���p3u��z�׿�>W�Xt�{�f���u_�:��/`���-��U$��z���ؖ���?�տ�׹�q����;5Fh�w��A��R��&D�D����σ.��dT����d��*U7�{{��L6����5g���� �"�`��C�z��s������eB�d�W9_jzSr�;WǪn?�qp)!�y��%\٦c��W�H����fV�}��i�kxy����:�iҰ��x������Ej�A���k�oI��_�Ƈ�դI�;\Q����I!H��J pwa���^/���h9N�h��r� n	����ȴ�<�yz2,%"��� L�<���(#�-`����ҋ70U'���ܻ�fs_��g�)�0����5�T��/O�����?j?{�pq�ak���b� ��";o�ґ�������Y�����ۤ�<Se�f�Ӗ��@g��*�wR� ���+��	�.X�u��"����~.��l9�LH���[�s���Kݦ�,�V#�����RkdM�u�f*�E79��hǕ�]HU�Hy�<ض�8eGv�q�I��U���B��x�J�А�bvGgI���C61�1��d(��*X����跘�Y\O�H�����fF�	�m�g䠐�!^��wm��=����������E8`��z$ުJrGCn��W�09����������M�
�5�H��~���/�er ���
Z�S���\'!���}��`��D�n_֣27g�&P�o���kF����\��5?�6�iI�G�n �� /���	�����"��W�;;��J�����g=����e�x0���Z����o�5�}�촌K�C���A�����2iƏ|���@��U��ꑔ��p���E6:ũc�e-�ʋ��Ĺ:{�=������(��~Ń!�kq	/UT�=�7O������U����^�����
�d�!��x�݆���T��b�!L" �L�8�զ{��ս����v?$�����/8Ȃ>�f��	���&b ���C����s�r� �C��M�?�-�B|���گ\�no��8�� ��;���5��oH7��f�n�_D��W� �0��f={9r����V����D��\0	{L�iG7��K�Eq�^������������[!W�ѧ[����4����|�Ц)o/�A|Vn�}*/����u�7��{zO����Õ �,.?�D2��'���!q��;���B�&z��}��_VL�}��c���(����(w�V�0�@I!�X��2� �-����<eR�-}��e�Ƣh|?V�{1���
������I@۟D���Y
9DW��f?&��*A��lƛ�(1_����!���U�ɵ�vL埍���$����V+'w�.�n��'�$3�Pd��o�K�$�44FrgF�n��V2�½`˛zqv� �V��X"�|��p�p�����=Ş%,�'���t�m�l��4��J���׳5�_�Dչ%c ���rH���g�>{��Bc�x�]��u�b���?ݐ���n´�L��f�ƿ�^H0���֩NLE�y��4W~��ö�[��i�M{�V��k��8����!�q��h��<�3w4��˞�Ts��k��T����~@��$-E@����2#7~<gKl��;j���n���8���� {��~�����ft�T
�����LOs�l�iC�#����p����+�Aͫ��-IP`a��G</�iUc�d;�P޶d<��{/�V<��5q�W�FИ�y�H��~X�K�O�~�0�'�:��W�t�|ხ#��k�����\��4�.E�4n�x6�QH�t[s�5"���ß6�P?&�	�ҧ�t��	Q��6[��-TґD[�v��k�ufV{�j�;�\��q�����K@#Z;䍚��	-�-~�9�j��d�e����OЮ�i�&�𨾸��1�SI!�a��g��p�ς�D:2:/�d�E�4AѬ��f�Pqq���s�O���l��'8ě�5\ߡm�O|�^�������"�S�8��Է��ْE`�������=��>%D
R�4"�	�.�	a��=AAmN޻t]�@���=�p�z%0Z��Hm��*����܂�W�Qj�K՝h�o�xL�� hqи3[���Yf�Z@�e����٪E�����7N�M��LT�	GBT8�t��(Gt�Q��&D�d���p�� ��J�=��V�?_���(Q����)�)����Qz&%���`�Ս��Z�TW���"ۙ�Җ���� �0����d�������(ԋJ�͛ch$�oG:ˎ�|�6V�+7�g�,X�ޥ���%x$���a�V/>����[�4�T��ᖄS�K�W�0§�<�A�L4���ɉ�Z��j��f�d��w��d��+�~��J6޿{~y�ԃ���d"�!��Z�O�짆���
d2��ޥ :HKb�U�%6I.?�J*�H�7�7/G!�2�AE��������܅P��gpc=�&c3|��a�K�M������
�6�|�Ȕ�C���%�/��\ˡ�����
�
լQ��y�Q���|�Bg`�,�P.�8݌�-���i�Q���7�R���ap�q�̵M�[ �w'옫�H����d��-�Xp6""�¤�� P��{{�����k�5/��]ܤ#j�V�m�"e	�	c謐���<�
ݏ[��8��(�W�7�|�����H~20�.�*EE��9=��R���s�=�rh`dE�dR�j���n��&��C	c6�_L�d���c/"	t����Qn�r���,Kp�گ�h���|��"D��C[k�]���d ��o���ߣ��� �{5pN���
h�2[>�]��~%x��&Nr�;�jF�ClN�i��30�d�����a��u���Y�f���*���BZ�+x=7S<��2� N�7ϺM�Xㅽ���cC������/o7����Hb~,�XT��0���2�FnC(��"���j�t���bW���'g�Z���e�Up�I �@c���[t.dn��̓)���\�k�y�i5��c���(�3-�<�&�����V�𖅉.�yK����س5`(W���yE��J �U�:&=��|��$�f����#'���;,ņgp%�̜�;�UU��e�'��/����$���_���nk4����}��p��I,;��M`L�r����铱8�nL,�\	��<��B�.�	?ɋ�gaMdv���޸?e=����$x�y��a���P0���7s�b�2���\�%t(mt cjP����u͹iR�k��l���""u��l>_Ȍy��rA�g�j���T8�{H�ih�"�&�J�G�Z5�5��B�ZEseDᤴ3�#�^��ތ��)<�!_��2���*F�����pe�+S�����V-G�t�j2�Tt�|���*��x.a� �J1�|�~�EI�wW&YUiFR�"���������[�z�|�;j��:�x��xn�F�{��Jm`�J;Ky�f����J�1��i/ZX�F�'�W���0"���,]w�\w��a��-��#2ݭ��vCU:To�p��G���	{���q7�iHQ����q�iMC?�s����P�\N����������5�PPzb,V��z�`�4�q#�g����#uf�;=u�����@�ET��!1�b��y�Я��B&����ƣ��С�F����|����O�v�����L����y{�)W���V�4�葥��ŰW�U��|�̳���{�����{�C�lF���@1�4����S���5Q�r*���O?v���c����["��(���@�ҝ�[ʶ�_?C�
j@�h!+�<��x��e4+{���� |���il����k�]�Fɑl�3+K#��J�ŔS���6��"T~�x��r"��	Ơ����*��)c#��d�gJ�*�8��|<�E�˶��ͥ�ƓW�W{�^���I}]:�Ʌ�/��ˎ!��]����2�#ԓ�F)e�_�6�Gh@�Zt�6u��Ϋ�{v:(eR r�+焯�"
M����l�����	@��8��#%��6�+LCKW��V M`�������-�z]ϯ*��%n��|q��\[�=�����:��Q��pr��B��ޕ ��S"�TE�Ɨ H�B���-�{m���(0m��qDB�5���O*(� 0Pl�I5xN�$� B/4V̪��|�BSkL/�/��F�g�]-7� ��dFI떵?Q�ߝ��,k u�-�3!�yc|�;v�l�1K�s�Ӭ�W�g��$@\2$>�@�1����8ed�;&K�%�1�`��tV�u�+<E�w�{�i�Z� �����-T�n&����p�L�/�e#��|�n���jQté�+�q��ľ6��j|�\�����xx��\�#m^}��O{fz��&G�q*���f�7����ϼ�uKf��_9�*Ю��(Jy�t����ik[�:7��:���u�ϸoE����|a��)���(�r��`.%�썹-�wA\$V��u$� U�>��Ñ�Iܡ�D��ص�t5��Be̥R����rG�D���C�F�}��:�h����	���2H|�"��x���/sX�����A�F�B@	S/½p��F���~�!�ߙJC�u�w�A��nϚC.�b~����;��K�wq�2~wop5:����^2o��$ȗp+�@�����a`D*,X��'��^B�xK��E��/�E37��j�6��*�� �fW�hB��8ϫ��0��N��l���+
��c3��w��LkT���� ���1��8��c�������WO�;�^��� X mq	�*�(���4��K<�%1��^v�����Ⱥ�Ͼ
���A�Pɦb�rZU�C|}*D'��x����Ma󋶸���cƭ[��^k#Ț����ƚ{�j�0�C%DV4���7�V��d�s�M\
���a��Q��-�XW����.�+dw7�P�����OLf\�c���5�0��l��*wt�|&�{D�,�{���x������ڿ;�6�~��9��6�h�2ڻK5���LV��p,Đ6ഭ����=���*��{mz�D�9�AwT�d��8OI���O��������F�W�VH��`��]s�`����堻�D�p���>&V���>�,w�E�xIZ��V8�ƚ�4b��۞�Oz|61�6(8���s����x<_��`j��tW���e��Djb�p���Ė r��u���7z�#S�7U�U������#��8 ��B��Et�8��R<�%"o|G�w&��YSEs�W+|�Zc�x�8h�T����������sP�X��b\�l��P�i/6��["����-�^ly�?��"�~_�����h2e�&ak�����n������J�gm�������c2�B��ȉ���>4A`M�e|���b���P�=!.�.�Q�ę����>��O&��s1|�^���/�j��x�����1(�/���8��w߈舒����s�Ɍ4gm4t]A�.�k'J���;��R!�u>��c_?L;��;��D̻{�ύKBG�2����'� 6v�yT��k����Uɘݓr�2������Bؖ'	+�0rߜ��*ޡ�����w���f�[̈́����ɲ�6�-����o�m ��a��\F2��dC��������؝��.RLŘf�\�F��V�Iv.�Co F�&n-S��2$_��K�0�$�OUą`�>�ix�j���UK���Պ������~P�<�-�zuS�N�"���)�g�}�=x2ř��XY������l�(��z��l��қ�FQhJk!�}7#sk�-+/v�n�u�����1��/���24�l@`%@�����x����x4��s�XY���-��M�-������L����x]�.O�e����W�H���d'�0O���a,�z㪷��nj"0��FWK��|���b�U�]p��7H����9Z�����"#���r�&�t9���*r�r�c,�X0�Z�i��x��K%��zP�[��;��Ru�Kv�Y�	�"��`�̔�-��|1-���C۹�_�5�An�
���H̩����CN����>�ۊ?�Nj��)a��TЮ(R�PLє8�|~���1f��8#��9��3$����_���>�v����D;��k3v����LjY��`@�Z���۷}/��_Ad�>�w�߸{�׫(s&��%�==>��d@8Բ�0�T�w{q���A��̺qa�Q����);l����a���RM���.�AęU34���9W2s�:�eW^S6ti��@?�E��N��Lu�,'�l%Pʹ3����+�� ���/|��Hl�p4pH6��P
Lz���N90�G���c+��p�2������Xuַ�����[]�b#����F׹�Z�]㼺Գ�-�/4�8��xm�MaXow��GZ������v�r�v�1�{�'H}���d¡R}��#�s���}�Y~�Ⱦ�^^DZ OPF8h	��b�\��Y������w�>e�!��aemd<�8�#���d9H�WΞ�h��N�˥J���,T�DL��}v$�̊�F2rk����]��yÑHi�D�U�;+�0�ޗmAب��'�E��Ŧ�=k�ë-Q�����P�m��փP��� �B������k�j���g�ހ�34&��Vz�F�Y�߉np�h�x�����_��К<���>���L�)�o������p5�9,R�t2���"m��cz�]�-�<k��>:���{'�M�kcW|CLfގ�|=U��׶c����T��+��.y�lV�O���g��/��rn�yd��o�t�{.��}h���QK�n^E�Rc��F���$ѣ�O�A�s��)��1�
�����P7�\��\�(��)!�U��9������(m��{H�r�	t�]ԏ���8ވ܉ON�a�?]��q}�L�����J�k14^9�ZSi��2^���8�}~U�ڶokF�_{F�If �\�ʾ�M��8R� D�3cÅh�	�>݀.3e`�6�;��Sh��Ӄ�����Tz��?�\���h�*"�$H"��	w�t|�K�x �{q��c�*��J(��2�_�z[W	 m}���X�hil���8�#�hPu���7��ձ�����ш=c�U	D�f����p���w�lvI�0�ʺ.�:�k���c��j�1F�N�2f���a4^<���Q'�	����X����lkAPziA��T��0����Uhc$�I���۠�Ő�ma3�0x���]L9�~��	�3��-��Q���e$������YdX���V������$�kĻ�^C�+u�?>p�&�� r����@��`r�"�DXm]ү����g%ó�x�>!}␏A���r��Wc#��Oo����;4� I�������Еc�Y������[�s��JR�XU>$�:����ۛ���wQ�$��'�6Ϊ?[ٙ��ͩj�������c�zB��N��s��\[F��r����S�����~~��$P��+�:잰�V��;�D�̳�|1;�;�Vʋ�f�j
M��Jq���W�DE�5,��������6��R� ��� ��?7F0fR. /�eq,�{�eHlT�Wj�����DC�<�)6W}Jhj�KK�קF,˭4���tI7~�v�$�GN�yn�%�^Fl�_Ve��v���9�^H�0���j8���o��9�x�Q�޹���J���R¸d�$��hA�����]S�-K�������B�]�J���A���/;C�G�xcΙ������&�ˮ)�c��SJ��C�orc⚼�B������D�M)�#����Ow�L�
0� ��Z�fo���J�x�t���q�{Rmu�L����(�_,������=����k���� �>6a��*�Wֵ�_)��\@�� �|��� ?��AN�U����C}�h�K�VCp���y�� �����L�\�\}�]����P�2����N���e2j��B��I��~v�hO��������cr�;�`4������v����#aG���U �#y7)W��U	#�&��RW�7N[Fo}{#���5d�IZ�Ft��!�����4�!�BBaZ�yA���V���`�co؆[r;�$�s����z�鶸�e��џ��q?~�^߰+�=��15?]�V�� ��7��x��7�������Q&.̰�����O�B�����=���y�54�wa��3����0���n>����볿/�t�sC'3�Br
<��:�,�y�1��r�Th�2ݻ���e�d�Ǯd]I;�J��J���W]d�"��Ќa�Q�{tX��a`���H�9�����! l\e�=�{�NP�zG��&�J�����o�O�D3O��f���[H�Q�3�*>�;h28?o�]/g>�9��Mx_�m%iTɒ5?�f��Hi2�E:�^Uϑ�r��R�nQ&��pS[(�kօ{'^�YL�@���F׏�B�!��ISrʙ7�@��z���c�	#��tӊ"��IeC|�z�^Ɂ�t�,����m���E���Z�V n'Y�e?�^c�
�d����'R+���)o�����{ J�����#�~�6#C�F�UBu�"}lQ���\"R+�Q�2����1�;M��X��a�ݚ]�,s��`�������ƽ(�k�i�m�Zgy<R	̦�&P�vC���4��V�Ja��"3�ٴ��0|=RX�/6Þǋ͍ޜ�~�6N4�*��P���M��_u�+�X�{�pi^}c �
zW1Ue�©F�G���/q��-��qp�EpرolA�)�k�`җ�b#
��rg(X���D�7?n1��/�\�:�7�Ć<�ÑJ�a������7�!Іy�q�!��*yN�.��j�.���U통w:��!£a�a�i�"�-k�D���+ϒI��ｶ�	ʍEp�5�W�E��:�V��XGj 	t#7D�
R��.ǥB�k秮QK�,%
�5\k����_3&7�����Q�"�Q�s��47j���3E�0uh�}k�6��/���R(���䇸k~���1��H���l��*VGk޳�.�f�hrl� $.��u#��K�����m�3O�O�6Ōh4쀌�F����|�hkJ��Ox����SN�XoW��sK˞���Űi�FeM��BG^@������!�ڸ$������>ׁ�(9)�@	<X*�0=X����������6�cz��\%+��6��6�^\!���@Mu�z6�M I1,�S޷�-�?��u�R�OJh@s����:O�ڊ�U���}#܎5�no%��3t�Ƀ)�pE(�f�O~�Zj�c�5�%x�
m���Š�\��
�6����nӫ�8�Ԯ1j/����ȃ�cˊǫ�M2�������c˛Yfq�+�⑺*˯!���V%e0�Q��>e!���;[}��Z����Ty��I*IE��_� m7.<N\�G�ڀ�b�#  �yc=��*idQ)i�K����p)� �6�qÍQ- [�����.���Uӫ�'��%.��Ct�`�q×�Z������WW�V��hÙ� ���� �ϧ߾<d#����1A*N~��j~7b%1�JH'�J`�-9���� vh���$�����c��l�/��wq׶��[k; I��-&Ll ����2�x�R-�������ou���+k���� n����vy�Q�s����ys�ՆLÄ��"UD�Qh�\��m��sK{��3H�E��_�c.�wF>y�we�-�M�u�p@&������-�%?4�B�m���2�$X�S޸���덳~��d+ȕrN�j��9�%�'6	3�������a�ի�a	���@)g��}y.�[>2��ϕpm����4Rd��)�He�^0��)UȪ������4؟5��4}�e������9"|SH9�2�
��EW��L�i-usZ�M�{β�=�;e�e�$��N����Z��~"�s�vVE�_��k���YL��|&SOƔ�r��'*�ODYZD���	sT��[}�����8��oz�H�6��M�w��������<��X�c>��j�w��pHg����N*��X�E���1j�&��O=�d +�� 7(j{F��NP���V.�J�%��JG�%�̡�R#�F�� �#��!� ڧV�O�)�8Ӳ�EcnG+�+��)�*��eS'�_#��V+?�Ha��
m�����ӥ�=�0��k��M�!e�XZ�iA5A缘V�����^�p��ҕ���G״�8ײP�9�A���\�qt?�VHo�� �R���$c7�C�o+$���Ӥ�o`q͓$��F�ZWQ?<�T��P��$C���ɯ_w��8Z;~���M>�Fg@�u�Z������*��������Q�2$�]����§�X�A�w� �����E�u�
F��Ϲ2��8�/�+��{��*q�o����^9�ܳ%��������jU�����\^"��ׁ�:����=�^���$a`�7	g�A/nC�O�L�u�����!I��7;d�H��_�l��D@�m���sc�d(8)�9���D����'0p�^&�_�wi��3���N��F��(��vC���(G��y�_k�S�Ȟ�X�1�~Ԍ��y����=�F�	d(�r�c���6�G���"~�36����y��%��J���r�-^DH���J�`
2@���6=�n.��y�\e^y�d#�D`=�fA��&�d��1��a���߳b.��.�)~�P�]"y�oo�xMv�MҜ4�<n��R���(1u�U�R?�'v��9,ў�p}LW*��2����
��I ���x�/����h�643���m0^FXL�-������J8ie�)wU�H�]�ep��ԗ�7��J����,hM�=*��c�vhK�~}wQy�h�������?HO_)g=���������� ��B��$2u+>��J�ޜ6�X?.�.\6R䅮���E���oFvB�rt«�]䈣�ש_82v��7��5I�h�=Kt5{:�_r�8m�'\���B��8U��W?�;���|M²���� 4+_�	���A~���������	G�A�.���T��}��H��UTĪ"/}4�'��#��F�mg�Gdz��G�.Z$W_)����)�BB&���GZYڰ�o7Ҍ�
�Iн�E�W���LL�*�1>T:���z���;�LHMs<#��C���_������JH� U.HX�$��O������A!B;��s�r�H�K��)O m���B-��!�?����q���V���B>P��!�`��XQ��'߅��d§]D	��|�dr:3Ml1�Ô�v���A�c�S��+G��UA$��t�O��q������2�
ڜ�Z��]:���~��[�:4B~')�r��Y���3��!�\���'u��=%*�#�~�>ߖĖ�)o���� g{��,dtɣ�C���	�������RF6�m���ؔ��R��za.��`��Z\P������p�� [�������r��0E�j��m�&�q�Lp�]=:��J��pG�ǒ�d	'/���R8��tx�{,�
���dYL�Յ��@T�5k��$u��'��GQ�o�c�d��L��Nr�'M�=���C��c@��1�w�<i�B�l�u�B���mG�^�:�YEt	P������E)���e|���
����n>��|��|�S���&q��W�nSG7�"n���4�T�����!���|�#���ۚPc���r�C|�!��+������uu:k��p��T�1����T||�{]�h�M� E	�3qyDx�(��[��r:.M��6qk�(&@�ۇ1���moW��z�(я.��o^���}^'�Vc�ܙk*�����@�'�f��#�ad�
O!/�"�pͤ��3Ӌ��L�`�B�3�t>���u�xN9,��^��9��{4��ɟ}�(U�����K}���e\�}�%���ܛ)��v����"�q��2O��V%`\Ք9�%��wBv/�U�^O�2�5�2���*��x���k�9�c�1-�Fc'����8��ٔ�1K��\��k��خ��0{`�q�x���Ie�#�1?�����oWk�f"��H����_�(�E�v?�H����q'e
+�wu�`��Yl��)$*�Z���Q�$+��*��`��s4|Vz6]&����c����HLzYSnH�]6:R�y�z3Y�sᖱF)�c��yT�y��F��JE�|	'�b���e��./ȼS)OX���k��o�x%D�-h��+u��9=Cx
	��rģ����-�y�G�␘GX��7�j��v[�Vo�j���ЈH��-`Hڡ:�+��#�����"֌�5�v�f���h�`�e��F�L�/�����	��ʖ*��L�@��ɑ��4-�[/:� ����gq^܃"zi��R�wb��ӭ9��TjA�K�q�w?�:�V�?�--�gr�w/�qv��p���`�9zf�hc;�Ф�
�l@A�-�FhA�Ȝ��9�r[y��6`����G��p,�͵۲[��1O��-5����M�_��ms���f.�$pHs�Y�$�pR���r���;�a����-�l[�Y`�Vk�܉�|��������-���7�&$u���I �JDL�N�w|K��Z��]��;�Տ"�e���@�'a��n�=���\q�պk�f\	� �[�A6t l��~�>ܝ\�ʉ�y[ڪ�uD��/wX��.pÌ��b��&�g����k��?�#��@�%���u�k�7V�����QY"ړ�L-��/_Sևy�5GS=�x��a;Eo�\N5���#)��-T��#h�۴�V�h
��xb��b,�~_���!4N>�M�E'N@�lr��^���[Gw�nU��_:�I�h�k٭�)����=%�?�(�����L$�Y|Y�%v�H��R����"������%؄J�Q6�wh=������.�|2zGa�3]�W6s�S�)!�/��09JC�b�V�5m�;P��Zܪ�����}���i��꼅���J ~ёv@ہA�S����P��yX5����C�鎭+��e|�[�!%:�SJ��W��i7Ȍ��Ȫ�F���'�-����j]Q4�֑��Q��L�R�*�~��n��Ak����m794���E;ڃ@��gVGB|_�e�-k��H�=��#����MK�Gb�[�<��R�{�vq�?��8�bL�{l�o4��"����M���L�;�Z-CNL�E���07�@��a������W���C>:�Jmv: $m�{�ȶj'����� Jίϟ��#>� d�dyW���0K��N�"��	�fm�\�Cφb褌�� �B��얹�cM����M�î����H�U���_��Ǥ�!x%b����AX��T9N�6�������kKz�JuE�)J7Ĭ��~ �\�f��Yl�睠}�4�o�к$k(c������[��./#u�'�d��E�2*H�&.Q<<��������2~���H���[|�. K+�EOƍC�2��`D_�tG���u�53�0~�a#���zbr�zz�2����%��&�z�5#��V]y0q���"��{�t���!1���Ƀ��$pׇ$��W��@�mS��-�e��Qn�fўsX��ъ�"^!I:���aߢ��<��H�	}Gv2�����)"��;�C�1�W�toso��Q"�hgI?
7�g�HG�D�&@�^\n":%Y��L�\-����R�W���o�.�5#��U���'ZeU�q,(�¨�kO0�0�-ON���ǵAe��P���[�AI��L|���m����E�k��w�li�;�>�6N� ��ZP��Y��UٝR�F��g����u��l�J�oH��|��t���R��<g�bw�e{U�h�P�]�gT.RY��J�`���Lx�~]���)+6A}�����]V{�WiS�:�=�-�P�[���p�*/�V�}�K���pg=[��
�t��1p�-��b$�Ȋ���:��1t E�EýI�b�SVL�c�eҠ�e���0��Q+9��� �!��8���?z��W@�V��tsJ����s��Lk��U/N��u����U�����n�m�N9e�t�d=J�yƥ[���u��Y��+@����㨸�^��3SݖN}����x���S$?q�,����mז��!aȺ�G�K�X�7�Yą�*zk�h��QVՂ�N/����a��Wը*��o"���30l<�o%^�G��%l���@X�|�!�x��9��Zz��ܕq���Y�㿎������,��6�c�Ҁb���$�6ۢh��ګAt��,��������[��0�'C�X1Π���&2
>�y�dM�%`�//�5޳�rFf��qƖbۼUx�S����t�����Vss�@��j����#6���H*K�c��,ݨ��mD�������:�H�W����ݪ��L}��>2a��2��B%����y�$��:e���y+cR�m��f[�A��t���|��<SBJ�7�ʤs����Jgj����>��qG�{Wdv��T���^!��f��Z� Z����B�����ʹ�4�=z��9�u�(�68����_FW�U::Tؤ`��8̤��(��TKEi�CA	�T�=^_ލR����ie�V|"�_���e�X����zk��'���V�CJE������^r9!�;�НN2D�"4q�KW�Ǫu�^��XF�q1n��T����싉{G)��!�͈@o��,hP|��� 
�7�l=	\�m��v�wJQ�'Dl��{4 ;Z+Aj����(���=rg��7��U�8�Xu��׫�iC��/@\��	�b�
B�>ހN�P�J_�<��`3��!=f����z��r٥�Q%2C���D�7�e񄦬{o3��z\���K��M���m�3�X	BΤ&Q��R�s�j�m�������n�,�� 
eG�?�xX}_��sG}�۫&X�.���=׼%��K�:\�^=?\��P����Y�k;�'Ƃ������(���s�o'���:90��Ak֏U_�""C�N�����_��8�K~^�5`!�9�@G��R���}^�S\%QK�|S�.��'9�Q��@HS鏞!ȃ�{��է�')@8��hk�6�#���Kɷ�WV&^�O���E��q��QC��P�L�x[��e���E���mwZ�S�A�2�H+7����N�|$Һ����n�ەkfC��gâL�5U[������e<�Ϳ��imD�D2�bcV�r"��MqRW��| U������z�L)�坦�pp�+Y���{��S�� %_��^���Ü��A��x%�ˈ[%n1�Y�����j�� ��;��lsr�Ƙ� y�v��&q��AOc�2?����3bʧ}*/^Y����t]�.��6MwU_fg�Yy����_�Jy$���������p� �������ٹd��y�n{�=�`J��N�Ў^�w���<[�wh�M�a�I	��i%t�yrp�)���>��ƛ�د�΁�{�MJ�4�(}�x�n��N=ˈ���B݀��-�Bnf�ܲ)�Z���Q�8�)[�C$�&<��Vw�K���TYk1d��`[R���{�bB��_�n��z�g`��jӺ���؏���e$��mB�;0��y�8Ɂ��!�B?�,'�s2�yV���'�� ۃ��.C�ǢôA��:@�8�>g����M���B�	:�pMF�7���uS�t��h�T��7\�a�����?�=Z��㶬�0T~��i,�=��Xv�sF����Y�H�F��RE�y��>@	�|1���SY[�t�V��3�D�=)$�<A��ó�d���������0��@M�Y�-_��:��AC��U�LL5�Y K�k������o�yK���Fs�%�zD��5_ڔn��_)�'����*W`��	&�了�>�'���0J�O��C���H��"$?�s=�ё����֟����Oj���y�hJc�%2��wS8�ٶ�#�3��\��
(� 1D��^��qZ^�k5齇8(�<��
	Ѯ�Vؘ2p�Q(n��k���|�tvsk���=eU6��B%��}�ik$׋���қU�y�Nw�i^G��}���qVQ�5��/2�V�p&_4�ղ#����r�}�[�#�0o�5�Z7�����w�lQ��DL2�L��f5�;��h��P�p�!�]n�I�V���N��e��O���^O��l�����H���+R>���1�O��g>�#��^�?�h�D��'����q�O!P��Q�E��۰nd?'�1p=`���0,U�Ij�]��_hj�B�_Bxg+ts-W\��+F�oHIu��m
�+0UrT�7�d�92��*�1f�?	���e�n���ڀ߻���4|� |� y���\]�D�W����O���Wԣ��G������=�؝r��g�-W���f��ܦ���Krb�����ȋK�S�ا���fIr�W���x/�M���O��u!��hM.� ���T�B6?���j �&����y��f��U`�b6�h7ča�K�J��I�w�An�Os�,Ƚ�uǷD���7t���J��˛45�������c��H".�WT�2U���6�b�V�xFڶ�FM�a[��_*��	�Rr��s.Mʣ��f�z�6��dle��Oy�gA�.����F�_	"���گ�I�1T�f���r���0 �\��˯�\�_�"Ir��{U2�x<G�!8�����84�U{ȡ�<~F��TD_�w^��33^r�գ�Q��r�O*�Qpa��M_�]��ƣ#o���Z~�ӛ�Z��t�ߋ�]�0H�>������J�_F�`�L�%�_�!�~�d[6�%+LXO��Эo�$n���`�c�:����'h��%T��>��4� D��I���e�t�K\��^�巀}Nr�"���%@������ԑ�������R�.�)��M��f�~N�s�w�OUv+��\8]��^����G�O.
���@����F"u��V��&79>N#f�>v�ުU���e��Z6�M��_��Q��s�h�1n��f�k����h��?�6�ڧ�K&,�9�<��m)�є�[�KK�/g��cT�bȗ�RT�`�����{LM�Y჻o���L�\�{x����t���(e�yq	N��R�=�0U���1I*B�)�<p�t�@�r2�`� C�tr#�g�����A6��U�L���t��!��TA�"�,f��s4A˃��ӎ�T�����ovdf��d m3t�i�J�3�O�8���.���P�Yg+��Z�k��&uZ0�9�eҝQ�����f4��,	U�$Q�-�n�y�l�!}5��:W�.�5����; �����q����6(&�����
`H-f�����@e�fO�a�����{/�7�~�0O0�8�P��~{� o�hZ����J��F_B�'p�*��FZ:���uL&54��긒����+�����X��N��:F�D�\�� ��!/��QOo_�����:G���sZ�K`cE��	���R�-~@LyĚx����H���Ϛ���o���؂�Sh �B|7"lp��4Vu��ϧ�aQ#(�V`ˍ����X��p��d^�t��N�geW>"�=��h�!�P�}����^�lFv|Hʪ�5��l2�]f�l�s�6�HP��6uo(� �m�4�u�̀6����� ���Q7ĕa��E�g6PM�r��4��/j�(%�ҷ8����8����X6��p�21!�A��d]}/�&����`�ae��GJ2�o��q����{����7W���g�嗖��Hs�X���U�0 ??S����xx��r��9 �G6Cw�b����P�kr�U����ʂ�ڷ��(���G�F�3Ӄ�omO�N����]6�q���¢k�F1M��n5�]��)���v̄#v�UWΟٕ�(�+u���? X���Zi�_��d!Aw��E�3�)NpX�$�����3c��z<���J�M���'�&'�vI����� ��Rg��z>;^짵�^��J�TD�P�ҝ���j���eeܓ�J}��fɠ��˼�W�&��V[�P���e�� E0��닸qd��8����N��Sj
�k�	��B�ϊ��s�g�NDL4U�,����Dq���ۺ&z)��d}�st,��{��$K�	H>���\�Ti�|{�����Y�'��K5<����b��&�)P��8�
�m�5�P�
2��~h��1f�{xΠȅJ ��i�2NT�
È�aR�}��@���i�T�L��^w�A2�[Ē�7�aIQW����o\B���-����A�wz��v5�es�>H{[%�X��!f�\ʻ�}�A�}Y�	Î�	�b��1w����g�@��|�z��mI�_��R�&!���*��9j��gy���ā���o�#.�d��)�o~���Q�_Bm�5),DH���bWZ+����,����C���.��F�d��y_;�����u�I܁���be��b>�d�R�o���[���'l��L�O8p$�ol1���/�}�]L7ǙLqߊ*}^N�r��\�&��,*1ɺ���2���`N��(����o�o �zh��3�DG�܃�h�{nGX�wz|b�2��a����X�3/�B肫����o�7�Z�\�5bZ��*����wO��{isFO����Dה� S�)>L���y+�W��-�RY�W��f�^�a>ˬR�78vD����BuW|�Z"���Pe#y���#:�$v��yE�S��~s���`䰓��B�7?}ͩR�N����9�V�nu.)��KұV[谢�n��dVGb#&�W��������D]@��%z�##UTK�Z����JJm	���3�M��k�a!� ��2�s�1�sXzQ�͢4�f���(�1H���0�T���g�+%��Bʒ���Rm-��e�����i[P�:�?@��8��=�a#V�B��<��6l�pƤ���)}�:ሐ+ݾ�feZ����uS�H��Q��3pUj�(#~�L�n�Q8�#9M�f�|����M
y��B�g��be��c������;�x,v��L	�(wQ�#�]���5RBh���k4��%m�\��n����J�����L9ϔ-���XT	S+�>�7w�H�k��7�_�(���x|y�=�w!_����.d�'F~�-�}D�kj��̇o�\ u�H��������С?��ř�L:ަo�Z�&ￍT'D	��!�tc����S��?+>m���:���?jؽu�1���*Mܣ)LOM�Y"3��v2$@	��w�����9�ݸ��<>���ٯ9*��e��Õ�t��m���#K�#�1ζ}<�t&`��`�.�E�W<y[2�[ g���)�f��X�
�c�~T�i����\��3,]elZG����(3��?p{���{����<��7���E9�_9��@iK���)$}T4�"BIZ5����Ԭ�%�Fst�(y�Pt�� �.���Ù����2�"�'v�<� �����8%�u��C\l�������@��JכKW��4Ԟ\:ʕ[oN:DG����3�*���#Jڧ�>���E�����v��M�`�lo���Jo�M�e2��m��ތ�o�nw�u�5E�����岣J�7y U��%rڲ��z���<S���ۼ)�&��n]x$�qmĆ �F�I�F����r -��-�A�T��;��=��}�(X*^#��,�u�w�[�q�Tbi���OG^�0	k�g0/�i�B��8v��#_�0Z��
�X#�Q`y����,�@к�����E���-8��2(F�<���pO���L
��GD�>ms'��� �{s�^��A\���9r9�w-��Q_���/0�E'�:���W�'�UQ����Iev���h�q��G�m�+I�k��\Z*UKI��7����Pf}�?Gcӄ,�){<t@�h�9�r#��0QJ\�=C2Ae�Z5rdA�A��<L�����F$�c;p$�ĕH�9q�Rٴ��t?*u 4�Tdq�����Ҹs~ʗ
�����
Yu���ճ�C�h[Db1���x\I�$<q8j�v�G��6&��9� ҷi�u�!����ie�Dh���VZU��[���r7$AL�G�ԀkCf=�*�r�>�3ˋ�!q��*�7!7���4>���9"�*�Y?�_#(P���oV�:z��x��]ebH�?W������)d&q��^I/KRu�A�[�n��%��v/ 4��C6��L�ߩ�кh��g#�R��+q�*��^xE��1������C<�;���Y?���p�N�
l�M��\���_tyXhG�u�o��s��*�>���l^U�	6�ⷫ�w�\�N�dŦ��Ph�ݏ������Ib+k�0G8��h��Lg�.(���y<�v�(���L֨B]����v3E�̎�o��r�p�@_��0!n�P�=%6��C�������¶퓝��}��T���E�_��1��������E�o����d��~��&�0���J��f��'l�����{�ui�h������`%]��3!֎��;
�&
�c��Y���� �N�S�IP��\�1�j�돻�-�RP�,PP���C��Ԍ���ҕ�K��[g#&fgʒ�ᝀKl0I&�{%d�p�>��/W܃�x&�LR'wS�֢:4�mJ�ns ���F��z��N��ܯ��C{,�ٗE]��*in�/2��l��R��*�7D�B�;-��@��Z�x#�ln�m,�h�E�u�Wd������ѝ9��á�Mf�D]/����|P#�9�4�C��2(N�1���+�Μ>��Nv4��k�0���,Sf�Ė�EXA��B�PKLZ�Xg��G6�������}��X���LݻG��|cH����=C�!� �_H��㐇���g�4NrQ`���:��Z9����If0��]ƅ�:*r�*Yc����n��Ѯ��X��3.>�$����b���M+�O�(w�"�d+��f�����%O4����9�������	��+�(�� E��u���{&�n���F��M�W T ���.i��M��=Q"2n�>�	�3ޛO��m�^a��}�.O�催 v��/0\~���/����h�tF�-��#ZKmMb�"�e�S�O'rJ �M��|��ǖ�h���D��6M���+,�i��\ԇ���&a��-��t��y�3����QC�M�Qp7J@bD��4:
�������Г-�Q��iDR������[���ް>TP�v���ӒJ��T���|{����Ô�PB�����]�p�R�$h���FN7<�=�7�љ��Ys(%�pK��	K�?c�I0R�xx�R���m����#�p�vf�FXD9�������~�3i#�ʦ��.��w#T��x��������Ƃ�Á͚��9ʩ>�f�c��iu������f� �2:�U|+���E����2_��z?Rz��4u��w�8��5~?�5P;�G�ݹ��#�+����4�����Dl8#C
���m��gj�H'W�V�lT���.�tTi#��yZ��]���rF �e��s ��ֶC`A�{^���-�ֲ�͏������Yn}R��X��kሰ�E7�r>�/���'P������.�<�
'��]������A�E�g�܉��w~�a$��b.G0�U8_b2L��hٱJԺ�GV��0"R��'L�e�!������FLm��=Y����bh��]W�r�sC-EW�b`Z
��X�Z��s�' XGD�B>l(�bqma�zM��ٲx4z���J�,���;����X��?q/�~�!�c��$}Z{ [/���O/��`>��/�<��dw��jyU��|����
�p����DT�(ʐQ\��և���mJV2�>l~�O*%����u��
�wi�O��׹��d�� ��Ϧ?��bc���I���w�����Mzq�@A��y�-�"N�u�Dx�K#u�ox�/}��(�a�Y#F�9�aj��Q3�ᬜ���]&�)�J)��2������s�}ܫ�N�W5�����)�j��$NwF�=���/�o��݀Kc���
�V˯�[���;ҝ;��1J<&�����jW�":"i[yΧL�×u/����31g��R�V���$��u<�I}��Ob�4�� ],�����佪��
�'�����V9
�|{?%Ъ?�6F�|9��n��Ap�x8���XZ�(�n��c��/^�n��t��2c-���^�Q�/S]�T�M�4
�\BǊ�0�����8�8��ōɟ%X����X�ng]B4�[vl�������/�.��ݦ�-��U��ZE#i���/"�X�.Ϋ�Q4W2��^�8 �-�?0�(�0����T�|�T0�x�LQ�;�S`r���Y=�?�'F��xի:Ώ]���[���k&5��̯��n�Έ)�{'�F�(�a��%��1��d������I#�m���8���!�J/.�(ܼ��y��܃{�i���}�!�Vg�k��V�v'�o�h�af�K��2&�ۋ���{�s�ݻ��R�vo�rz�]h�����{v�_�	��@qd4�4�6�����]�L �N{!l��9��h�kgQw���H���AH6����:��`��
:��j��$�b���X�jR�K� ����xF��1I6H3h�5���O�X),�>;ϳ�ꫛ������vDy�Ij���L�T�2�ӏ���F��66���?4M�vƮ^v��'}��ώ��\�n�-���tT������,�~�A���Q�)]*�E�<ጞ��ZO[S"ߍ
h�PU(�D+��ޭ�V\���&5�?Y��RHM�M𮅓aHHͣ�l�V�!Xa�=��c>�WS-�#�M�
b�ˢ����?,o�����&/�g�( C��s"�B�V�:IU5��Wo*8���v�m*�l����,�(��j!�B;H��	�3�A��,Z.�˧e7�W}rXF�U8��+��x��|��BF[0�:&�S��<*�j�=j(�J!z�0vz��k�4o���q��0��%�d`�c�
$v��r��|N<�rK.��h�;.d�@ItĚ����Z{-�~�o��Y\�_��9[���F����c: ֔!��L�M<�����[�fF$a�F-hK��o��a�c�09�Y,L˩t�Hc��U4׬x���Mi��B��ta�!�M�yc��B�.V���'��+� �B�O�)`=�XA]4����aT<����4@6�����ae^2�g��e޾�6�0
	�PS)�L�s5���+ƺ/�u��xRgz"��K���f.y�fi�5�_ 6�r����}s:(e�Wl̃�1�Cfs�>�*��._���i��=�><�Q�����h�`! �m�c/染���r �˾9�@!���LE���`�^���CY�3�u�J_tg�V�$�y< W��bҭdBL�DYb�A�?fe�w`��f�RK�1o#G���Rٍ��a�2����v���ǫ��؏��๽�'�-�d��'���7j�[Q ?}����/���t�IK������4Zgv��7�;��s�0p{f�y����![��������B[��Zf�I�Δ?��3�gT[�d���n�
��p�:�@��Y��-*!�ӵn�R��*3�kM��(�[���Ҍv�a��<�dGD����ds]`���5��HR`7�s9?�ƛa��Ȧv�$T���;U���
<͙�(�T#�TB��d��\�  ��8j��}�&�͓�
&P����/���/�B�C�ge{�2�;�I��ש�U��|�S����1E��b�lΜ���8��8��Z(*�8�2*�yI�ö���� ��D�)X�"��D�OrߐS��5�Ǐ�����|��O2x�c^���5e�b�� �b�}8����@�[����~���j��.J�/�K	����.���%�ePl��^��v�v��8�$+o#��%)��?`�2�10 ���
TX��j�_�1HB`b0�?h����|1�q�!�WY�3U�W�?��PCn��g�6��i���w���U���V[pL\��\x��6j�)2�1�X�)qF���"�'K�Lj��46�#=�����I
��B/@��]��<!o�d�^�Ť�Z��7�B�f�,r�W�hN;Q�v��߀�v;��"L�`��t���r�:@f|��&�����L0�jq�k�`9��c��mA���b��	�ʔ�I��_5b����1���흦7�[w���v���k]��G(o7����oޥ�ֱ��Z!Kn�:U�p��)��V���ʯ�X�&�=-��+�����Ͳ��l�|x�jH�����q�i�G�>>6g�ȴ�X6#�	"��������k����+��%�T��j����&�J���$��mB�(�ə��bȔ?*A���%�l�}r��ؽ�ƴ$�stV���r���\�.�Ę�aE-�}��߃�\�����_����(��w�(`��a�ї7����#��h��"�T�?�9�ʠP�S�s'���T#�����Ng��`�O`@Yt���������3/No�� iQ�E��� jv�!;|��%�����`d���*����c�8wV4�����=����X`,�0g�y����X۬��L���:�I�����^6h�GF��	�C�%�� �9�J|+
�PL�b:��P��&�Ue��6\����I���s��]��e�LRhz◕�~w�I�h��Qv���)�Z·���t�k>�_������owsF�}�Mhv�%��Ȱ��J����T����)̤&�������.����^���(���.�C��wA�^�Ԋ�bfO9�_E�$����)O�*"w�Q�5����v��b	�=k��ʓD�w\�!��Ȧj#X�8Ո�t��-�l'���gH���cٶ��O�|���ƞ�<�S�D��-�@�&�d�Z����e&ۉ���Ֆ�:ʹF۲�W7q��[-�.-LrF��^Z���a�)�pr����a�9��>�<�4�F)�⯚�\��I*�%ќ5���˫��̀���_�u� ����K����2��9�LӚ���0s|�L��1`��g����ƃ��C���WPԹ�>l�d�n}c�5��C ؛����7[�E-��\��خV4p�3Ǳ2
�G�����`�ȍ�6�p_+
��FM �t��d���l�ݠ��G��f�)�� ����!r�%��T�"���z+�`�Ǐ$�"j�w�`��Ս��r�{�Z?<��V��(�^����F'�f�B��u�7����%� _)��ϱ��L�`����P�`��i �#�o�Z��gI�S����=�F�Љtўm���=�4~��k�@	�m���u�kJ{��BF���s5���CT��c� P=��������L�)(.u��X�g	�?�y>��'�q�wU�SU�Jɍ{���3D���b"������۽�hY�k=ԧ�@��wx`"cb�V�L��'��`(�d��E`YN�����X'N@�	td賧i⊮,���r�=p���9��/O�
��<ŀ��3���������d��7��M
�����Ur�2�d$�lq��4�eԼ1�؃~@ �BDh� ��	c����"�)�t��P(�*����a���/�P�2QF1:>��d�Ή��}O��i�UUƽI��R�"� c��?A�(V���~A�`�p�߇�EJ�o� w"�rr�CAB���ؾ�� �����|~d����y�F��^k#k;��|��Y!p��i�ֳ��ċ������W�KM�	��9�}aG!���D:�}%0Ի"�����z@����2f�+��iS�&��*������l��n�F�s�p<�5�����
�����}�����5-��ZnNe(#e���|��V���<��+KE�i\V(j�v�E��e��+@Q��#B��)>��6�q��,06f[-�V�8Go���l;���`]���3l�$��H��6��O���Pm�46�R8��m��4Z��LD�7 J~�L�R�wmu%-��z����z��n�!V �HLҾRJ(F��8��ZQ�,�4��lz>m�m� ����x/��m~�JͮxG����'���i)T�K��df����X��� ܋B���JC���4
��a�;M*���B�0D�����5L����uͽ�06�����=�r���K����9�5� \F^�6�d��#���LH5N:���^���ڕ6E��ρ�s��b؟��O�|�����Y�؊r�jX���f\/I�R(|��^T�H:º��S/�����p�	 lB>8|�Ea��D���w�h�y�G"���}��@���mj���>mVt�#u�P2�e#֙[aCO|RD����Pߕ�R:�IKE�\C�ߣ�{���I��`h7���S��� R����Q�IđO4(���\�N�t�}�_ى���1���u\1�I��`e�!0�gku���Q@(�P��:h��d��lZ>���fZ#]�$���?9h��a�`���Z )������U�< ��S�	Gq9�X��}����ݴ��3��2NZ�����	܈	���i�GK���E� ��P�{W��SK�mң�mc���Ų���.�h�TY͔b�:��S1M��#���L�ҥJ�(�{(��R� DJd%��ڕg˒uΌB;>�����6�*�_� Du��F�?�T���}+���Gg�v��n�1S_V!�D3���7��"�U��:\Gi0�ńҹ���w�>v��@���޸�O��"����#�,���5��"%�5mz�톛Rq���wN�:��"�K�ɩ�\?7ƕX�uTSB]������A,z�U���׭�O�Ua)�3��[l礿%��PS�\�I�;����QA!0'n�m�[=�\U@�{����s��C�G��P�
����k�y�G�j��s�R���!�������Bmլ"_ʱ��:Ɲx�j| c���F��6�2�e�CKŊi�2Z�M�p����CN>�����`]�I��c[�����o���XА� IV	�IU�R���uZ�&�~�S�:�:��L|D	X>�߈:�6�m�f8!�p��ipW��L��[T�҂;��t���#<ؤ���OR��$:_}��jϬ<��(�))Q*苿,Y����f�������8��	�Lg��]w u�16��� �z�����3�}���^���4�Oҽ�{ok��4�ݐ�[�� ��'6'�bj>�e���a�rˬ��n;X��:ߌK�B�ق��B��V�[���p�jX�5�`u<��#m�D��KL�կâ�����ޗ�y�Q��t���|Gc \4F:ʜ?�Fhip?�4�i<EU�&��x+@?����i��t|�:�7��]�jO���v�����ߧ�:�Q�G�/I�@������.�iB�����(�X���p�����Ɓ(��DVQC)[��ʱT��
C8�19*�((����|y��QV'u���4�<��3��B�g��z�0�f0���1���iw�����>+M4����a`�yh�$c���:�����'�vp"�bs7� ��̳r׷�*|���{S<��>�(��ɷ07���3@(�`��6�R����[�-uy;x޼HۘBĉ�NgV���I�09�4_�O�m5Z���6!�%��"�
90��/@T�'ô��u\�%s?��w$.�g�~���0xϑT����4�!�`�Ł����#���k����t�o�f��f�x��H������\�$2ez\BhrI;��J+f `�WꉇL��xL���A<���`�,�#k/,�	�q�K�"�&����j|F" ��I#����ajB�S��m��і\�?�5��_�2���oH{���JACB���-��:a`�7����y�e�ӿ��}�6����Y�B<|k�� �F�)���9̫���\>��+�jgUks#�����[b/뽧?�Ab�� �0E�S &!�*��]s��� B~��X�'v��a���>q]����J��T�������ؠ���)Kg��C�w���Sh��8���s8s:;��o�OB��q����#Bm#��qU�L�Z���a�.>I��� 4M���p��v�~�oxi�L��L���#\]䄡�c6u2��;�K�󁨓tc��w@�O��`;�'�Ch��0Z�+��2�7��D�� �C�UE���݂�m+p�O&���V�t�e b�dZȁ1sGY��m�j�ߒY����K2�9�Gްfrn���{ �������Ժ823�^R3+Ŏ���������Tϴ�ч�H�nx^�u/�M�eJ�_���yV`�v�ڭ Egh8�k\�i�xR ��	g [l"��M	�d�I �&KV�c��W��~�ϝ&��
N���������_�$�ϴ��{Y�c�fOQ�.�/�/���*��@J	ߌf9��8ۈ}�zf�kS!���((�������jjR��KW��$�:>���hd`����T�VVv��EsÒ?��"�4��˒��"�j>"��/��G����h�		ه�dMf�ꎓ#/;(onψ�J�C>�ʄ�n"Ǹ`�=���.�}pnZQ>2��p��)*~�B�/�;_�ǫg�:Ϣ�G���ta �]/�`�������ş�1M�OF�e�"��n��]=,b v��Q�u��22
c�j�����dfUF�L�]V���~��%���8��κ�lZB�����=Rq��<Oj��)�}�Wyr:g��0�� h
^R�(�~��8�LnI���Ǉ9�U�W��$�1�#"0,�Ħs1��7L�,���Q!PT��`��@,�a�:�xTP#oCC5���t�*_U�]"�t�A�j�\���-�K1$q¬Cp�Q��	A ӱޯ�|������!��$�^:�QO�J�:�C3>����u�D��*�a�	A��[<^��P{��� ,}4�=�W�5g�Σ��;��ߕ�؍fZzF�+���<����Rur���v�,&�J�kfcL[�6>�%#�/s�������K�r�Ŀ��fZ��쒶lv@�P��̯���p��%[����0.^�<�̵���J�;�D�ǲ�*҉�y�x�1P����e��M���+��mD9.+�m�荿�<��R� 6l�S�P�9.r9,Ø�7��\p�O����2E((�zU��d�9�����.y��U8Fz��lh��h�?`��h(?�D��o����6��_A��V��A�5�z�4�5GԐ}���5����u�u$��u�-�ᾎ7�g�( l � �=$���T��U��Wm�����<�P������߶�$Rwt�pG�"���	���zi �2���Z���z)iΒC�xu�dN6�|�R�&캳J �5���(�U��.q��
��	,!����k�Ƭ���6�:��kx�%!o�t�Z��W��_�/�V�V�E,���쬤]9(zmsX�ݴ�\t����3O�u�:�ÂEӽߤ>� ���֑R��p��R���
��#��=�����>])*y;�#>��Υ����=Ry���5U~첻�O��wr��P`91���T=X���6������_{Ђ/��%6���(������l�-��R��`��3d��_�L8�|��󕇓��.�I�f��6��ӗ��įzv`�I�>�D���ov�:��\�~�:��%�
�'lZ�#�'}w4���`Ȳ4M���r[Ң���vL�|��?���ؑ9�"����c���n�'k\�E?
cz�Å�p�0u����o���4˒��W.:�6��8���.>IZӱ�t�lhOP���ܱ�B/�6��,�]�:�߷��]�V�:OS{��8��q�eKL��q�3�O,˕x�0D�1�y���EO/bDv�R�z�^�ew�E]�����gl�����gDŅ���0	��ԏ���G�`c��� �L�����1~�#�=���J<CM'���r��{�T1�6�	�S_�Rf|��ju���
�$�!���3a�h�Aa�r�&��"~=���N��N�&��	��,�)�>ꎘ��}I�j�/m�W/<�nt6��~�1�2����H
����Hs���E��䥫O�>LW�Y�l��j^��������b_ۭ��V�ƀDg�8�U�NS��x��>*o���p{���f@�����.\� �<n�[�N���
4ׇ��b�5���Ȃ�d~��&�	7��!�T���?�
h�O�
��z'9P���$u�����/^y��=�mpl��kg2��8�\�a�e7 �R�8�l8�����ӏ�rg��>y�^�pə:(H@5ڬ��5��II��i�${��6

q0�u�
�F*	��&c%���Mpĭp�^�LNՆ�d�|D�ό��g�&Q��0XX�}�NT8�c��9�� ����rN�>�B['De��ɿwK{�xȶ,]��R6���1���4k�3.��a�X1��a�C��2�Į�Ұ��6^�h�ɝ�\e9��3l�����9�.z�b*i�LĞ�'��Q�Q*KC����㫽��xrk���s��2�P�jࠓ���Ic��ak�̯�E�.8�����*���׍y�Ls�RQLu��<�l�,�!c�V!a���];�D�4����+�����ï��OpG����v����)' |P ���e��C	7ߢ���Iǁ�8�����RQ�ޔ�J��F�4Z��n>r�F�w�W�T����Fr�[,c��άR��W�LL�һ���g���L��V�(1���i�,*�2�KF�&"�)";�O=s��M�##�,R;���6St�����b�gµ���=���D���vO�+ (�'���:1������a9d�BN~%s��9KLS�x����sM�q���L]���EVÀHGO+�M%���j#�*�	������LS��,�/1�����T�C7[3c�|'	J��#ٮ�n�SAѺ�<�e���H����Q�t�txGCL�V��0j�'8&io|����r	U2:x�҂1��(Nh�؍�.��q/��܃�q��U��׃�T��pW́,S��:�0�U�`� xL�?`�D��IF_�*SN�>ܡ~ɷx�&V}Y�'i���*��HfF�A�Z����(�=�}��\�q��Ĩ��{�7���A�&\�WZ��O:���y��j�eS�/(t�1	'�(O4~>�Hy-y�j�ŋ_���W��b���t�/g�����YM�N��U�j�ˑ�P��l���I-�%���?K�x�[����Lr���g{jRӓą����z��cA�U���M|#,�{=4�Vh[!58�,p�#����4_&�ÄC�K���5g�4k��Ul��S��!�50�P��ʟ��{i�
7�Xp\�"y<���Ɍ��wo��p����qdZ
�t�?��)��3������8�qua!����͝�\]ğ`1-ۯ�c��F1s�Xm�I���k�u�N��s˵����,{����{0ܛ'?��y�B��8�#8�!�][� +���Ⱥ4t�R�I@�#�����XN�tO8mB��H���^O_﷕p}ס���c���U��d8��V��VJ!�!���F�"�RWc����iKH��,i��٭�ӓ��~��Bd�߁����f*��9���$��S���A2KsahR�Մ�DV�X��s�RMT�:x��k7����e��0/�Ɛ�ܟ�G��l#�i����F�e_%��2_���\Ыm��`�3�����JFˀꦍ�j��K��ca���M��G�^�lN�g�yu�E�^�	݂�J�����!�ݰWn.�OVw-�Э$�#K�J�V�d)"�F�jE�@��mJ�{�ND�ѡ9����Z7��ƉE]�y���8yO�\)i���ȭ�M{q�T��2�.	o.s��ω�����2hc!]�a�^����f�:���I��ۀS��_�i0��f}O��%8<ӛG����@���(�+��%��v	��i�'|�I-��04Uvdb�9���p'˳ɹ%`L�o�zQ���ѿ�1����Mh����:���Mi�S�k`���w�x�hݽ�J����2�	�`хl���r��W���,�L{��6C���PA�h��ӚNA��Ĝ%����A����5au��Nk�'�Ds�.RC*��������Ĉ�Ro:��:X���SAv׻�u�x��}A	�f����ʊ[b�0�¡.�R��� Z�WG'�bh�_����Tk�+�F�[���IH�vR�~�1��*� �z�=Ix󔈟\"�o�}�Vi��}9��s�$���^a�4cд�$Zh�Y�9�7k�M��D����b1m�/n%�A�w��6�,�3ܰЫ�i�ݭ؆�(HgH�㩯�͖� 3�A�>Aә��t�� ���Z6��5�����gړ���Y�]�P=�\l^}}�,��e�Co�X�Bs�ժ#}1��hnL�N
��HObd�mF���4�a�T$|�������M�Z�%_��(�����Dr�(��	5�#����B�:��7�pNFq^�o q���F�\~��]�)��!�p�C��o�`�SM5���Ŀu0ٌ���Ǻ�<Ȁ�Oi_l^�Kp��$���s$�J!����|����]�V�巌Ck��)'�|]�o��XX�b'�vk��tN���5��v����(֥�N��SN�w)b�w@Ҹ�YH�!C�L0�#	ȉ���!I�� $Z�=Gwi�<ߍc�6��k#{e&��~8ێ6Ws�jF�w�����^��a�uc��;�5�� |uݔv��풇���}�c�=	I�������,k���vQ�dm��~C��H�U�T�����ݨ�13_1~P�@���^��X�I����S3����7QF��V���2�kqZ�C��'�E�§:�Yʔ�Q�,Ü���mje����u���� ��ֳ�ˣ�?����fg^b�6��=>�\lJ�AP4|�&D�8j����r�J���eF�����g����(�y� ���L�u��<šo� ��)+ʕq�Ǟ��:u�+GÉ��j��Du��c��I��zQ�y�'��o�~K}u�9K�J�
�.�8��N�D3���8q�Z�t���;}Ii����Z��K�ꃯ2���s�5t�R� ��<�v\Z. xűO��x���B��3�p�r?r&�{�N��ڞ%:I�q���=|R�Y0��G%x�̏ZEB�V��m��-��Ԕ��?���W�{9�̌WD �����K�#�|���п|9a���Z�0�ɺ���)- V�&�.�
�&��2D��'qF���Ū��>�"d%�?a��Q���"p���\R&I�m�� &�� *�[��v�*��H��Ӷ��S#��%�l�~+$:."D�t�a�����C��@�D��QZw���I����0X�A�ˍ�e*s����i��=��v��&|S�<jL+V�h��V�Z�H���LL��>���V谤����I�~���Ut�6���$������z��}�l}��B�O�5�\	�V��,x��V})�8yo��ՠ�>��/l/�!�V���'���i���i�zΌߪ5 m1**���j����-Sb��J|l���<���\5�g�D��p�;V_�1����ٹ.�ޤ ,,�&G�2��!g	��yz�Ǝ#�}�P����QZ����OQ �N�(�[bVh��cJoA���*�`*����#���rל��£Rg2!�O����Cm,��'�.RP(�"�i-/���U�r_����b/Ip��u]�\�
y1�v�e�7{�-c\�����f�).�0�@�4���&d�[|"uy~T�Vd&l&��"`�ܻڐ��2Xh�3��A�YX%��PyM^�I����;���$�"���L��1M��uY%k;����u(��,� C�;;K3N�^l�kZ�;��"³��q��k0߹�w5޾{���T�%�Iv���g{@����ϼ�(@�o�g͑�rv�U���K���B�ω�R�o%� �Z�c�N���B���n�����ZK�}��|�h^���bƎv���S��K�KLQ��Ԝ-�Q�k������8&ihѰK����J���Ԯy�{@~��S��G	�̞��U�>riaK!R�B���U?\Gr~C[�*����~�`L�e>��ԣ����B�i���A�PF@:�b�r_�,=����&��Ч\gmW�6�0�AĿ��=��>�o2Aֲ>���𽎞�~�t寯��E�!0��$.}�<XΗC��Ka��`Ñ+Ғy8z���uw"�vRd�rD�)�O�ݾ�u�*�����9�Υ� �!�
r!���+M6�ߐ����6b�	2���ſ�@����p�9��6�S����ُS�sGjhѱ��̦0vF0�L��f��&�,`H6��$���B1o��/s{�&��	j�o�	Ss�R�,����N��F:5��l]+�m���9^�:��˄�m?��P�I��$���\37N��7�����A.q )� �.�ucw	ͦ<a����/��]����7�@r��}2�x����I�`#DCn܊�p�k=Ō�ҝ��c4�M�Qb�ӿ1��
g�zt����6>���ꄿ��s褄����W��J�oE�T�n,^��+��ɾIN���5����z����i]JVF�oH�p�5iS�z(�D���r�-Ȅ�("�G|�>\�g&)F�<���t�A���Й�!�F��a�p\�U�0;Ѩ8t�O�fk���L׃j z�_�����u�b�g��O[i����*JT�d[��_ɊR2y<j�<6<������iUX��
l7z�H-�W�j'�X�zg���w%�Ôp�T�)�\K�����0h^6��y�jZ��A\L4s�U
"�����f���3}��HR��n�w�}-��/��i��k�38����(��8v�:*�9n3y�͉�{�7�6��a��b\�Ǧ��+�Ql������[�ƿ�f	�q�4]�ٖJ���'T�X�lV�RhV����B�B���`w�01��Y�!L�F��B���C*��&Z�o��Zw�Ç6�0�������	�����y��13�DvG�b[*!�2�W?��l~�^=�,H3K�6����,p���~���t��ԲD����5f�E���\�ZMp��:ځ���\,*S���=���'�[�}�|(t�Ok�9)�\�q%<�S��ĳ��L\ɚ���bd#�>��bͣ���g�B�{!�4[C2I�ĺ���+�dv,��qq�p�1��K1:�p�L���O?�R{#�k�Kx�h�)8�GY
p����x8E��!]K6�V�r�Ta(z��8\�J�R)G�u�h�����z�\r~�=��^��'��s��3������x�~����/��g ���$jͽ�5~��tF�j�ǚ���hZ��yKG7��y׺�,P��_����]�}5�a���EN�m�5�aG1a��o�MTx\p��z�ҠX��PK�ӱ��L��I�P�/}��Z����ؕ
��R�����]h��[CWl>+�:�VQ�R� �1//4�����[V�o��O|�͡s<og�!l_Lr@��^��A�ka�F����6��'��D�>�D��Ƌҗ4��"�%A�c�ܠ#���bl�4�DTVX(*ݠۚH:�Z&��7�I2��Q< $��)����\wN_���T�����z����߈$��	%�ЂG�ߦ3��f����(�k<i�w7���eXj��WE�u��DVд<�9%NL\�)l]�B��9�./�C`�Uz&��T��0�����#yA�p��U�\�����Q���"�I�% |Q�Zf�g�"(���'V8�W\ %�/z��o���ќ$/@�7��.��̈�)�y������ϿKY�&���}:'��Cs�b�GP�C�����������<�b�ֽ�k�d�N�1wɆ�wH9Mh��q���XNM?�)�$0����;%��2����"K������� i����0���y]ǽ���;�tX[,��V���b�S~7��\�|������o����wBEr��+c���©}P��搒����wq�t����HM��Z*8
`��Ha�`D��W��`m�.$3�*2Ğ��>ͣ�ϕ�0���M���89�����L��"�=�ǰ�t=:k��3K�֙�H1�w7 �j�ʒ��ɭ��RF8�l�k�����H;�u�9��6�d�����֫�TA�)�$�B;L^��?�>z^,����cAs}z�T2�WxL�%��|
n�'}J���4f`�\�VL`�⧞���S�CŪ�&��[a���5 G{��O�Ž��I��+��"V9�(�#��������DzKբu����S$�i|�\�0��j�%��o�(n�YI�|7��0̕ԭ�au���\��B��لA���rL�L�SA!� M���i7*Q_a%�b�Tͺ�Jv��j��F3z�G?GB�֘�$����6@|�+CS�*�EC1��nU�o��(	��$s�2�U{2l�}J|�}D>0�W�b�XJ��ITd��D"9���M˞?ik3?��9�ְ&P�?�W�N�
�#7˻-��1��k*�� B����n���<a��!
��;@����I?<t��U%�|wz�ڪ�,�/�u�����-휯��ԯLG�
o��"�Z[�,\��-߈$;��6�?)W��+��@��
�Dx'֭�Hw�H|j���Ȳ��>V9��;#�GzAvQY~��=�ix�q��=ϧIƃg�p3�'��S��h`=a��{&�z��]FUTRq�l�Q�#�ۓ��Hp6�C���L�D��`Hz9#WNWO�Q��ם��*�(r��y,b��5�,�}�
�R0���ό�]R��+��$�0D.���j4z�K����U���L��ׯS�Y�r������o�|v�ƍ��n����C�UY�����%R��mNSi�V��;qu����BWK�3������e��ɥ>�&[��0�ǧ�U�3~@s�jM޸ڢRZ
3
��doyT�����2��#
����~�_�S:�~Q(�	8/�ʽ��@9�3��vԼ5K^(8�D�U1잝{P�;�܍�x���V1>?���EڨA��tľ�ͼ��XV���z �	��S�h�J?�{X�y���{�\M�V�oͪp��,}�X���-+�L>�������3�׶>���Z��+�+����o�8��#,���4��%j�wh��'ю/!k�&��?�;���&�d�[W�Y��n�M��Hx1�H�0�A6�ĳ;�]N����k����՞�ٴ�'Yo�~X�FG��>Ҟy|�3�q���0���y`��d������K��]Lp}�H����x�E��o��d7l��&�9*���*���In�q9j�l�^r�P�H�1��*+8p���΄�6݃��MO|0��%�bb��d�B)`�j�2�ۂG�B%��
(���0	��*�d�Fe���sEW�e��|���ȸ��a��Cy�����0Ӣ����d���e�J�F#Bl�'���;�H�X��
ү����ޢ+�J)m����;ӨJ�Zj\�~�e҂i
uaOV*U9��U(���8�CA��D���&x���NMs�b6�=��mV�#�Ju�TT��Я��1�?���D���r�p Q�D9:a��4u1��0�ש���?#�7?��
m_�Q8ruI�#����wb������G����d���!�?��Y�)ka)��xK�/��+4n�Ҕ���������uT=ѦK�DD��]7KZc�W�"F��ᅫ[���6;%h���# Tr,�fN�����f�?�pm7�o�U�j0��ɿ�e��~���� '����DWW�u��C�}�_�Ⱥ+�����H_TuX5�#)�A�43�f$˭������˥f��@"�� d�d��U[v�@}Q�){P,&���f�~��
�������	}=d(��C�j�h��Wj���@Fgq8�ܫ��T���bbM�^���E{Z�5 �;t�k��!*P6�e3�C)��s�C���E�/^x�D�����<�ה/�*tN�N�����휽�D(p�=��zr6��������d��ڄ�]!tsw��OK<:�袄w�:mj_^��|Zdau�7�O��fTƓ���Y�@ΐH'�f�*�*q� :Đ���3����B�~�Lp�"�d�)���g���ɬ���F
m��۩��HZ�E� ��A���jj�b��Ѱ+Lm�J\��~:��o	�!�[
���Sx�����!�Ȱk��2���Rz�
�'/�Vk	��� ����rh"�*�6V�[�6�f_���|��?^�W1�e���?�P:�+&�k�ՎT^ϳ��)�,"/0A�)Hĥ�˛�ʣ=u�5���a�ɗ�;�!�?	̈���Jd2<_�;5I\h" ��C�kA~��Q�E�	kH�U�UJ3��Ӑ a\^߲mO|�$U�A��>��s!�"�e0��o�,��Q]�N��
οO!��N.�v>�퓞���Ѿ�֮QȬ^>�na'}M��#���ᣞU~��oj�7��W����:.��!Ȅ��'uό�|�L�����Up7��A��I�7�bU(`�g.����L�?�B�kb��������>�d ]t�r(j?����`���$��/,��������	�.?�W�؋7�3������0��Ǿ��i�+ ���5`Y����0�+&Ϲ}��)*�T
��n!��n۷b>�0CA�>� ߆��H=�0����*��f�=���=�w-�0�����c���'[�qxD��I��{��OAk������Ǡ�S���Φ�kpf���V.Z8�*.#�Y�j�!�i�`S�fO�Eb��`ˤ�r[��^빑<d�5EYQuj�$���is�7�edz#s��c��z�
۲o����,A�jU�χD{Ş�49G��y�iP�n�����]�t9��/�u=�������仡ĭ���ЦR�;/����5��ٛ�����LL���U��w�7b#��)�9l1xVzc�&x��g`M'a��x6�8p� ���L�'�T�Ϥe;���g(x鯤e�ٓ&��L��2g	_]�c~r��	�Ws�?U�|?M�	B�͢gd���(2�	��Ĉ�י�U�.�𤿇u39��fEŴ?����8z|���Z����-�_N}��0{fŷ�6��#zkk�ܮ��J̟K�� ,V�� �����GYH}Xz\��զ�W�9;_�(!�ߏX���L�|���i�W�c*�}]��jp���H_�'��F)�C���@n�*�������[��ʤAɰ�:�l�w7��6��DRSǰ\��+�S����x�ƏrE�+b&	�0���k�k�OB{�61�X��}<����Z��=�P�zt�$x5�m�h\r�/u����e+J�H��'D�y��!A���Hј�3�۸��tE #5-�m�-xo6("�� W`��F����M���:�Q��2�C|TuN�{1��~����>�΂��@� �1O�g��(i!+ �{�ƔT��v��Xi��Q\�O�vx#�Ý��xfSa!`��]7�Cc�Ѭ(�X@�0�H��n���X�m)�':��~B���\�L�hY?|v�Ci��@~}$�J[���֓N�oޜ��%Q�">]���E����>n�רې&�͎RC�Y��t:��RY*��]b�@�Ќ�b	��z4��Ԗf�1��8��Z�@	�����\��/���7G�����^�t;L���%Ҋ66g��b�W#4��¾�����\�61f]���9�>:��e��5h����MzS������!��7%���ϭ��I=���`��M[5���R�?��L���ci=�i:�/�꓂1Ӳ���<&�lҺ!���c0:K�^�3dU��轜�&E0؀Un���ͩ��@�=�������/؍�OOLk��=��x�2V�>����H�����Z����9��تGM���1����d۠|qLb�wN���{���B�1n���G�:~����H,�0<(?_ﻷn�}ϵ���(�p���7ݎW��M6�}띅=�xT-����U%-�R��H%B9p(-.!�tb�a 5��TZ?��(*Z����c.�-qT^_���=��myͶ]�)y�,Y5��=Z�uYf�Qsw�[/D�c�f��S;�[I����yST͟Fأ�*�+��*w���X�Soa�c~�KM�:�l3sD�(��Z%����2x��(���q|p���̎����(U
p!���tk�cJ�_5^�o���F>;���f
�eQ�M<��bn.!���,t����i�9/��-��{0m0J����Xx�p�i3B=q/�6�ɫh�P����3}m�to�S�S>=:wM�����V#Έ{�
s�[
�e�JW.�`O�ePHSQ�a��&@�rkT�e�*���'��(��ћZ��gm�+�����R�1��8KH����}g��T����s��U?y���7�<%��"��r�ұ:�fk~�|��N���2�#�2)��/�k��6�J4�t@ޞa��E)�[L[�?�Pw�j�zU� k&�7�4��o� �P�/'��//G��<w�����*0H�#�@,bdQ��<y�?.�o�*�cߛ���)��:'\ӹ1��_ͫ�����`�`�RǢ�17$R8�ډ�˲*Nh�"���^����Dx?�f-��k
��ݫ�U��B�(�j�:qhN�0NN��H�'�4��aŋ>��?[��k�z�m���7o݁TweȵY�@�T�jR?��cG]�Y���D���x����:5Z��+3K/��c�^�����M�HA��?5�|!ld�a�gu�J�)L�/�Iu����_�$��0hZ�����Pn�/�w��c�gW�(C�.�����nE���!��JU�����#�8	�;��d[W�����*by�ч�{��qM��r��,bs�}�����we��S;��2�2��fL��%\}�h�(��,�7�������1�p���t����19*��M,r ֍_	3�*q\����A����puI)V�p"�O�+��ȉ�JO�ϛԾr�{	O*<//������� Xp���xGPW�h]y>Ҷk*G�ej�bxm*���-Qu
kMi ��	(H�n�Q���M�~����W�#z<������N�����g�M D��vj�J	����F+Hq�>�FHB�d���!�X6(a]��{���G5w4��:o6��^���2��}`��aP�[Rڛw����#�E�f��>�1r��	!|��#Z���,��dI�&�~�K��3�K���|��j�7D3	sq����H�����/cP����|<���j.]H�KO�k�:���d�o��80�� ]nm=��=	C�%R�
 e»�8CV��)�O4�P�~U�C�����0Ƨs0+�_��r�����ǚ��������N<�i-8ي���U���P����ĭ�W�~%�x[��8v�9���K�	|�8n�!�d���T8L.X���Jy$1��n����������ƹZL��b�����y[ǋ���}֟F�t�0���1g��^Fc��q׶
!�8~s��J��4TtQv��؄��cp��3��[l�l_�	uH�J��U�ӝU�zf�1����������3c�ns���ef�vJo+�yN�����(T�����`���X�~�G(@�ik�aLۣuR�EG�r�:�J�3�.ẗ́dVf��S��j��w��ت�� ����R�֖>z�lS m���~�U�`��R�b��d%K=�7�2WS�|=�	R�. �EE,��4�1�&TO|6�ѥ�W>:쒆�jx�"kI��W��KԱ�4be�[L�����G����D*���>��P�}�K��(�Д�Htih�I58���!-��KQ e2�= ��i��ؘ�z�%�Y�E:�Sr����+y��;�`t#����up�4�#��?B0i^�n����.�ZN��W@��n�Pf핫<v�/z����)��u	�H��F�g��e�a/��l9):y�/�á��R
�ӓb�����Ax�}b:�
y���+�6i���7A����w��:�,Rʷ��+�>�K�3l��|�'���֨�������!�(����%�i"�m�XMv��2�82��[É��K��� ���QV�$<�r�f��nH�D�>&XeRب����µK�/p�=���O�`�=w^��Z=������l�E��H��U��':�>�7�,�G���n&"��0�@J
s��	�BQd��N�9�N(��S�E�Fx[rQw��<�H\R�g���"�Cv'���\��t.,V��v���O<�UZ��6[|���<\;y<�\�i-l��!��,[�{"G�T�����'G��q�B����n��PJN;��
c��zF�d��и��5)쭹�b'�j�ըy�t �̔� ��wmW�Қ���YDn>�]��Ӹ�͐%]�(����hb��I��a�h��y
���F���`8.����W!a��*����!�6n��m�F�����)�Y4�EU��Yd�|���XC��]�!e�qbr�$�p]û&��ڃK���r��Mלk��)�?������. �?�Kqˇ��i>�b�S�)ʰН���
�C�n�\��/�^��Q{���DhE/�/�T��1�V���a���%u�uEBʻ�N�V�;�'Dr�e��r��ø<8�t����"ԑ��U(k|��#N�
�I�Ct>D|�l��w���6
��3��z[��DfƢ�ǡ�l�����6��yց�2��L����Kn_ k��XsT�@/h�<���4���m��TD�[}�. ���A��M=5U���7,�E��Cp1��|��^���hq���8p��Z�����+��8t�
HxF�\�*.BKE�|�����ȃ���D@� /�Q�X��*�j;�$.}N)T��4I���T�.��)�g�D�*����Gw��i��.*Ǥհ�mGK����l�����˼)Y.�b^�@A�<��0l>jfk��*6�ǒ��Ū�ԯvVկ~ψ�˒Yu0�Oкq�𷤦� �ύ=j��(�3���pg�s*�/�VG�A��؞p�|�eր��OK��+��Bs�Ȇ"f�-�\ɭ5����x{n�\���3Ȁ��{�%Ӵ�cj[�g�"觚�l����Z����>�˥P��M�dY�mŁ1��3<��u�q��Fn��qhy�w��y2`n�R��¼IԿ8C���!�Xex�w�Yj��fPK�\u��E�u������7��3�WD.�a�sRJ�?�x� �����?��-�W�-��zth��SS*�e�]~�{�3 o`lcB˕�m&�:P�>w����S�֫���z��<���`S�o�!uF���^V!za�U9�U�ĸ����}�ޠ3�p3b��EN$�~�X�žك���G�e���=��vDռ�Ǹ/�sS���T��-�+8S����Yy���{�Bj�݀�S�C�����wkzY?��т�5E�@@m�:��!`=�Bo�.=a(W�b�*FDz��񴔉Oӈ�ŀ��A�p�]��Ao-2cp��~'��T�n��Y�I�M<�
PnZ�w.����!Vr̸��9;�`�ϻ���2��^�/GL�
A-��_�g��.j�g������y�4�{�Pډ@A�u]j}<��'c��{Ձ�x�\�׻��c�&�����k�w�����<�[u�Έ77|���v���y����{�]o�N4����.Er�ޜ@$����q�ͤ�<�!�Q(Њ^W�܈�X��Xy���.ı����y��v���q;��*W\��)@��5��^E�Յ^��kZE��^�ՓҾB{L&�.g؇�0�6ϚS����
��5&�+f]!�#Q�y�>�x� ��� ��=Ū3&Ԁ��$|������2����AB���2��5pY�K�&�tϾy���
�}\]�@�S=�j���7Z�{
0ħ~2�!F��E����P�?���NDG�(ӂ�6��+���b�\[cT�f��h`t���KH��0�f�i��q��ͻc,��y��K�M1oa�f�k�(�s�Lj$������D�WK��sa(��̕׽UR����i��Ӹ� ��C#}ى�L��s�E�NRE���H���\�l4�^��Y���OĽ-z?�f����TǏ@Q��q4o���v	�uf��q�Z����h(�}+-*�*fY�bȶt�R��IF��[�B�N��N]�
�DKG�ǻ{E���h�q�s�|c�4�F�nRa�%�ko�󿳬ĺ��7F���D�̱q%�،�8'8��8A�%��+1��_\�D�!	�j�%դ��lF=xhc=�T���_8/oX-��Gq��T�"aA��G^L�ٍ��_p@�B��:���vFE��2ϐH+�?��$�zz��9�Ҍ�S�ۘ��t���9�q�j�5��7�
��K4E�φ����e��DY��u�Ŝ_轆ў�F�i���(b�RL���&�r��(�;F�n�t���1mҿ^���d��oh�����a}�w.Y�~l㱑yE�K���_u�&2Ă40�WWq�!�r�i�k��F�l�ء*���M (-u������ۀb/�6]���3{-���Њ���'� 2?�Uo�6�����rq���#kC��������]y�ͫ���Q Sb��0GuM�O�o�g��+�}�=wnBt1d�Խ�۶gC
�����bE�F%���2��~��*��-��|e��5��-M<�]wk t�V�h��*��]1#��I=`т~y?f̲��bn���8C���{�w��zٍAR�:W��͎�V�)�{���}b�-P��;,�=�����ʀ�sL� ��w�T���p�(��#*:-G.L�5-L��{S/�Ya�*��dB��|S��l#���-�OЕ�,>Lp $h�(�[��r��mW6�k�0�e��L�>�/��j������d�T��MF�x!��t��J`?�+�L]G?�!@��k��e| �I��X����$���B�~s`a��eT
KT���i������AmKR!�N,a���E��$�4��˝������r���C����ݟ8O���G�S�/R�-�,��7�i�&rQ�29zއ�WP���-s�o�ukJw7&���<�%O�������3�\$^����f�k��1&�q{d��,w]ꩻ�⁸��#+%��#8��b6���vk=�ô�uQ:���:0<w<���nׁ`�X$���J���!aj�Ȫ5.�F!ϫl��r�"t�T��-���A�,���P)����;�	�¹C @�G�����٭�	(wЮ�O���A���M`�I5�#'��3ۿ���]���q#�I��w�����7J��[;�����%~0���z)���^���@��\����-k~��1��յHf�<ip70H���gX����t�AH���.G�=Y��PQD��r#h���~2��ݗBe$K/�6���3�Ԉ���s�������ߝ5�����L� �N�;�=�Q��jJ�?�
�`5���j���nT�|�C;�Uq�ȥP���]�`��/�>�/�^�
�.����y���9"Mܛ([��W_�����N�.�i�@ӔO4�_�ù�+�}^�t�vpC�ۀ��(¾�-��!JD[Rx�1P"��(�*�
�@\K���Y��$Pު`N��|QT��G�W�+���ٰ�f��f�E>`oR��)4'�/yy;�r��o_��g~[�W���<�AC�?�J����R#�^����L����ў_'f��<%JL
��`�J�������O��`�XhK_P�% ��.%�n��b�۠ט�l3�-&m=q�����~S�,��k��Q�aL��8���`� >��Щ]�˯�� @�������%t�4VCt��j���˯8*^�Q�����n����s�ȣ�Mz(�2h*аFӗ��C.f��a��"�*)�D��p���q5yܱ��Ԓ��&!�<��E�\G�G \UO8ͮ�ﺶ��X�$@���Κ[|����i���pͰ�+�&U����ͅ�@�����Y`i�~�O!�B���0�\�s�l��'�`6�Mz �p�f���c&�&�=&[���^�����
{��N��N�p.�r3�&�!?O�c4��U�T������󠅆{I�e��	���%�=�$"C��[շ��P�:7�Dq���=�OY�#�el�5Z�]y:�Q�TM��D]l����/�@�8���j�!�]�����m��V�k�ww����>���يF0:�G/�+9匉׺���K'�S�h�=�d
�f1��}
��v��/K�4p4���mFX���x�1����B.���b��q��,V�d{=ҿH�`;m���4TA�(��ղ�j,�ɵ�:6�wK|� |��Nu4�FP��"�"���К�y+� fl���w�:ϗ^��T�(2�P_w�δcP2v2��#���C)�K�rE���1]G2���G����WefӫO*}9�r#NP}��-Y�}EW����'��TT�˲�Q$瑭]�2�0������� "���K����'�_hＵ�t]��p��zcן1�x�ZCU~I<tOR�ԡ)�v0���+�FK$���)ʌI[]��\G,ɹ�0LD�o��(\�u�_��ۓR̫�o��{��_���=Fq��d� ����Ք(J���e���q�A>���sM��dZ�#���%������o�j~�GquM�Jp9k&L�6+/ͳA@��WK�35�Z�D�p�i���yW58�f˞C�h?`�����R��Rn�Q�P[~���nYX��̉3����$����G���%m\ι/w8����g�� (�M⵰�dim���(� ��4r��κ[��	��~�׫��ξ�u�6U�G*n��(ۛf_��!Qj�O_���o+�dB<����B�V{�~�x�ϝ�4��`�)�>�zu$>�;]u&��O�kk�c��z� �p�������v���4.���Z����8�s�:b04�W�x�V�QAߡ�"}�'��\j�����T���H�	B�K>Azs�W]�E�D��r�C���Ë��9ү�P�Եڞ���"
n�w=KY�ڦi�2�ؾ�2�HM�s�'��E�l|�n_����d��0r��Y��z��W� ;#�R�,�[ �����i�*:"\;��in��\Ҧ��6|i���E%�^`��󣯾�֋a����lBA��g�{�4s����KD5������eh�Z9�ª�@�o�\������V�a�Zm���2�f���Z"K���E���D�;ɩ�@��}�%ra�WS�y"��"�"O[�K�ƹ�P�&~T����e���DoD��F��A\v,�pՃ���l.�8�&�#W�
�I���Y޷��#`;�W��x
Mֹ�/Z$m©�!��>ֲ�%�`*p��bذx\��`�1�n���'zf�/�,�U����T�v#a�+8R�J
h��|
d$S��8��d������fD�+���%�T�8�������Q��o�cI�_C�y���褈�w���T4#r�`�E
>k���[H����{|	�~-��ԋ�1bI&KBk~Mo�UY$?��Q��I(��m��.�Z��ѵO�!�]��n[�����d!|�0X2dK�ſ"a��v0�m�>5w+/�h*�o�Z��,t�7t�0ٰQ\+����0�[�$=�e�jg�-��Y����L��M���!���S@�0"�,Y1eX0Lc�VZ��0W:"��5��̢L���ֈ�/vO��.���HLn!�X��E��?�U�DJqsҙ��u�Id�N�?
I/�Fr�,��ۡI��a�<,�G�[nV���3a|��ҩ���ͷ���\���/���Ƽ㩸�~�Z:�#�8�8�S���������4�{����N�0�h��o�w�ϕ��7�&�j[����,c�
dT����O՘OXv���i�O�YC>���9`�2T Y2üT��\��n�;����eGf��^�����o9��'ܳ�(�ƃU�Z<^O&��	$�s^y����T����&A]i�t�ȹ]Ve�޻x�����C޻�3�����gQ���:��0i۲Jh���=��#p�^JW.?���������Q��p]��g�U�$���0�L +�}�D��[T�3֔��m$�-8�ě��W��W,S��ߠ��.��Y��L����C��5T�Tg|���-�P�5A0�@k��a(6���2�y�M�M�x��׫'-rE���)z�Õ+����@�vY�D�?Y���I�!l���&�<��S��T23��":_c"c�ʙ|`��+�C�4f*"V?�xMj�
�����g��F�i��H�7�v��D�FK�v���~����q�����5V&�Hk!��"��a4�Z�i5��G
Q�ě�1�EU�)�A�~HsN4G�`2��&���.� �3��Q�0�d��[�-��~`F['�r7��� u��sko�"y�n���P��=r����+���=u����&�x��լpT�ص}4�P�Dn�(��7�E�`�-� ph��%�;��䭨�Jߌ�<̭U�Z����h!�|�\k��b�f�zuY��z�/���Ŏ��)mn��x{�`�y������ݶZ{V,	F���DC������� K�ɪ$	I7|%:�U�?T{T���ln�N��F����Q�j�L��n���4�OrL�k@�O�Ѽec��(� m^ZP�L������-�.L�n��@y
 �In2=g��F���¾�'E��<���Ռܘ��:>�1���D01�G/���\�&�p�jp�l����Wc���b�or�S��
�K9�cT�+6D�ױ��7�9�B/���$h���|W�EW���zZ�A�3�{�6P+�h[S�`��z�_��Utt�y�w��/��oV�h)k��D&�$��1q���i����̮�lƙi�/9����i÷�p��IM'�Ȁ�
���zޒ�]s9�^�P*!/��Gut&��#mi���+��4|�Ի����
�ķ�`t����{��*�Iˬs��P�[��7&*���f��?}�t��' ^��Km�?d ?��5s1���\M����%}O�@�e
�VPʢD�ьP�̸$K��5+���Pģ32��+��ˑ���5���Ih���rsr�q�˅*�)�\�s�]8�bz2��ˣ}]JIiL-t�!��F�j@h-�j���Gd�?|�y��v�"p��c�͋��������fJ~��,Y�ˍT�%���+��}�{xE�0gQ!���*��f�s#=":�(�Q��Y�7V��Faļ]�.�=�>0�K}��ۇ��a@�K���I3E�d=aC�何��ϵFC�������1<�A�a�%_��4A����`
�E�ۖ���#�q#��o�x3%��<�����<�3�*l64тe�yH�BJ�����YUҁ����a4�	�"�����8	��6D�bm3�53��6ܔi�ʟ �֫/Su#7y��҅� �s�/���މ�SY�OxD������B���a��c�rǳ0:�S��ܓR��Ȉ���%k�ߩ&�(K��,�����"���d8[�fd_恞�&MeL�e{��qV�94;E��j�S���6���).��L�ʷ?�6�%�Y�~�Q��9��m��5����e���2x�БƂ��$.���[Z�k�O��@��H1 kR��<�R���)2tj��G�%UV�p�)�|`~��|l<ni�(&{������(���k��<��~�h�J�ɳTl��Ga�;+::�=Oh�$a�Ouq����#;�t����:,��:���ֱ��b�ԧ��D�jE���e�3�zX`��I�e��>�Qn���4#���wU�V���/q@��W��^u�rH����j-��:�sK��?>1�;�G�~n�í�Ƀ����	��PNxә|��Kr3��,ލ�0����HĽFCW��*��7���[���ŉ59�fCv.��L��5s6h�n�x���V�:Pu�,Q8� Le���M[ׁ'S��&�� t�B}.
�!^/kql9���z_)���+^h
'�HB"U`I{� S�W�����C"�w5��#V���9vlYQ�C/=)c���לx!!�%��+E�F���� aՌ�/F�0я��F�U��2�aa��:V�H$s����Db/�Q("���/"�n�0�s��D�A<n4��`��J�6���4&ZK �W���*󿂋�_��Qo��[�9��`�����L��x^��r..
��rpd�i��"����)���	8��L�oC`8m�6A�4n81^XY,g�
-c�/QR`ӕ�ʰ����_�}�Q)N�Fp��_J{��7��.}�QLc��߉�aD�W&/�Hl
��d�S|9������o.O��U�Q�x�Q6��g��ۧr��tpe�/���6���W@a{��{xäζi�Ƥ$;Us
�u S������o��Ih�6^=7���j3�o��d�m�8�L�y%J�%��j��-�r,&xd�-9����YX!r�Q��pC]��֧�8w����_�\s������l���֬bZQ}�����	J�c����>����ױn[��1WW�ⰲ�������)(r[*��sZ��<��k6��0Ю��@�Y1Fp��i��= m�li�@��,R��D'?iw��_l��]s�k����J���o�;ԋ!n�4{���P�Ȧc�si�S���6)!#�x��X�����VF���f<��4��!�qF��
�m���A�m�	2+��Ґ�+�c � 9{kx� ��y~��wٽ�h�$���8J��3	�y��~�p��<��5��|�>1Zv���Q�<�,��zf���;�Վ=��!�%n���Z�V�@>�%��{�X����*C�L���kж�-u���僈;`�%-M/g�W�xUOy=���^�V�VX�ov���<�ޘ�����n��)��jC�P�g�?�>�G��[�.WC�}V(���sBn<�b(��$�y&��)V���-qV���M�+y���"Qxa�H�H"G��V�o�LA}L�x�ߑ��;Q��EˎZ$����e�]�gy*Ɗ��T�f�1���Fhĺ���V@a�������}ps�B(��{�>����j,������"c�Ls�����<����xb٩���lg�7�.��m?����8��!�8J�8��C���������1;�����2�'_����V�Ί�g�����'b5b�T+�40LH�x� ���u���
�(!T�y�ų���0��(�,��6��aj���~�$�~�I�'����܄v��W�����I$��l� ���AI~�;�ȃ�j�;5��2�T�;�Y�I-'�3IuJrՏ��uO�@�5�����xc����tp�����n�����8����k�P�p�[����*�jA����r&�
��릝�2�T����c�'k`������Ԙ�±���1Q:�^�q�v����d�Q ��x�>�6U&ԣF��v�0;�a���lk���d3Q�&�^0k�O-���eI�|��έ�o��߁;LE�Y ��l��i��
n�i�Y<�m��Bh5�RG�ȍ
_~顛��G�X�'��TN����|���,1�]��o 6�c)���iSa�?�d㩸���H�F�����oo��X_P6�T`nKx��'�mt1h�" �̷i�;5���N��@�f�`�כ�н��;��x6K � ̣�����h��3�����O>E�Y�rK�D��P�h�"�gl� Ⱒ���~ ��� ̀���
���l��_���Yܗ�ɤ��on�T3�"�@\��K��������n�k���Ρ1!��jn|� �n�N��09,��S;�00��_Z�3��9c��m=����6�b�(y{�5��_V����-�M�4`��kj�?�_�՗��4	Q��k�o�%��OʽKfi�H^D6kڨfKy��$���Y�/�H�ؾ�!�U��@aY�.��:�y���V~UIs�ځ� S:��T��H&{A�o�
���y��7����SI�O�"�XLMF5�)v�Lr/����i(���"��О��O�f����9�~�EA>7#�x)��� ��꿷v�[�ǯ�I)�%<�\�:ܖ"��l�s��NS"䅉_�յ�ˀ'RKἂ�W���g m/����������A��_������On���:�թ��E�.L�i)�[���1­�4�x������h52"/"����c�&���E���l�"�Dx4������Ȳ���q��P��� ��G��8��^O67A�F]�B����d������Kտ��(?�)*Nϡf��zGR����w�̓�]�4չyIZg��x��ֆ��]=�3&����'j(�ޗq���ޜq���Ϣ��t��7 ��OȐ$�4�S@�G�5�F���
~��R3�@�,̕r�PȪ��k7#��i<I�QPEC��_�u��!)Y-�6���* ����_ӷ�F�Ǩ��m�g[��mx�~tZ��IS@Vɥ3�b]~:��ͼgo���A"3W�؊]ws@�OtlM�T'��lf�,�/��~�����&�Wj���8�_�[
�!�-����ؤUs������N�Y❋��s�R2�)����~1"	&n�*�Fn��w��������yQ��M}W3 �(h���" ~��sK��LZ'��H=d�Q3s[�r�5��]����E^n(==]���O�u��g���)<x�
�AO�&{��yf��R�R�n�b<(��̭�$S�GC�'�2o�F������M�%��)�I_v e*��O�ɷ����x����Z��� X��;�����VD��= /]����F�x�2o�L�y{���7��/���#C�8q���e<>�y霡���	�B���V^�{.N�	�U�����cj8��8|�j	C{�6��r�>T!�&4��׬̉�Z�ubl�H�5��T�Hs����Չ�����h��4�#�9_Bx�:F� ph�`�~s�K�Hjt,��\@n����_�Щ��a�GղA��M�d8�K��џ�1 ��*?<6��9���C���7�k��>=o�8<����-G��yϢ��O�Ur΍J0z7U�]jpG+|f �!{�`��)��NB磖�7�yY����gd�`����� ��p��f��5���o�j�G�j��\eݷ��С&8T9�S"����3�hn�Z>�~��.�S�`���Q`E7bm=|8s.u~��=ڲ�k6#�j�7ج�nI��_���:�t�f�v�p~at��_�]�+��$� �I��<ڽ�S�!���if�+�0}.�_'`�����0z���J���{�Y8��ûpA{�z��;o��"e|� �vCs|LA�ibd�q�b��z��.�ۦ6�ޛnW���[�^L�?�e �F`��_������1T����
�����Ė�kZ:���
P%��.#�Q4)雽�
I�̻~���+�s�D�>O!>�����؆�|�2��T����'&����L����� �o
��"W�Ѕ�=\��-���É��I<��f�v-;�2���.2��=hzgVS�>-}�Z�kI.m�p>��ٷ),�R�H2��?I����d�~n0w�.p����?9%��{����Bi�jud ��q�b~��76��XvPu�2����wB�=����Y'j�4���X�������d@T�G嘦.��3�2&xN����=�/�c�4-X�O������R���np�Q��|ke��1�H�)�~�-���|��Qd}0���5�!b���@�2��ܷMp釴�Ș�ʇT:�_�UBW;9؟E5V8��/�O0ex�L����>��WZ�U?oأV�~��Q[LѴ���w��Kb�nqQ���P� @���E[���5V��C��Z��V��ȶ[r=*е+�!/t�[�wE�?�{�.�p��4�,0��M/�dÉ�6�ҕ8�w����2s��zL?��vT/��f��]��>YH)�m�ʥJ�d�l8�\�z��_Ct㪝���m����q�#R�a����w���и��wKh!X�!A�٤4HX0	�Y�,M��J�K� /-ġP���6־�$�|�L�TC� H�c���p#���6�oԜS#�2VR`wF6�0�&��
���06�ؖ�r�c>�}�`�#������k��,���c�LE��,[��E�(��5�f�(x1�� �q�e]]�&�3ۯ��`{2喕�����:��j['��૓l��պZn��I�WY�Z?�5���Klʒ����Ws�n��aM�SAc�R�*�_Y�"Gd�^��y�Ez�[y�ȣ��pE�@�pC޺+)����} ��7z�U�������q���� �v	�����W��і��fXn
�LX=�C�_���\ˏn��s��e��?�B�=�����I�`�Ph-��w'�}�-EҖ��!F{쑀;jk<;��r�L���7�2��_��4W�T=�����&����ΤF���]���WEu�Ǖ=]a�!l�L��qB�Wɍ�S_;*r)�W`�P��*5˻���H���bF�[�ܲ����)�mB������ݛ�����D�^pӡ�O�G�)4�P�,�'�V��N����|Q�x��df�����޹'�2"��{��U�*�_�Jy�b�\��R���*�!oؕ(�����8K�}j�ׅÊ�o���t%ʯ66,�F9Ns��c��X�oe��%�?� WN]\a�.�H���n�W3c�
�+�@��: ���ه�|�Fsf�B	Ng��^OeN��&����<�e �|�_ �kgu�0��/s�s��t3��0����l�o
�G�.-�+�aA3A�\���� *��*W9�>\V�}�b���J���,���~h8z���^�,	7��AD*�5�<�vJ枰��=Q�|t�l�Z��R�~�~4�"|ڭ�a�З�9�{\�p�g��z��'���1ȃ!�ҼR�S�Ժx�U7��J{^KP��� �u#4��u�Iܡ��1����e��p�cu��4�@L]��`E�Eaiw]����N��mr�� ���,���ƛ�Hv�kQ�U���3A�^����p���ͧ����h"��쿺 �ZP�H��S�<V��U�UqM�Կ��e"�b�������J4�`�����t�?�*�tk�g�
�*��q�/�ȗV��u�7[e�+<ZV�s�!��ƛ���[�L�a+��}�pܑ���J2��Ii�ڐͩ���%��F��RBT���.��<���,]�O�ߏ���TrC7p�����t���G����7ka@p�i��"U��
����X�O�r�
�&�ء�qId�n߉�����e	+����a�lK�
�LK�qUH�P�6ɘ�c�j�)��)Ó�#���hq���A������7<1���=�4�`#"�?p�8�;
�A��%wMLg+.�y�
�����a=,�	��O�G�F��e,D �Vwi+��<{?P���!�ڐɂ�Z�;�`�bT	��ٹT��L݌����ses��K���΋���!�m�`��W������G[� ���p�t�*&��沴�y��v��O��-�G��4�����P <�(D_�������@NU�4ʻ���0M�f|KJ���)����@���ӭ���Ze	��-���P�E�n{���Y��:������gi�r�cO8,�ʜ���H+{��d�%�P�W�S�~o�H�+������.BN�#{7��Z�{�b:#03ۖ��\��f�c����ڋ�p-�`��<��N	"gM��/�y4Ov��x�[��(#8_�ٟg������*��ܵk�n�j��\�0^�>Y�����4�{"�N�dk���y[���&&���_/�[�+�(�yC����&߽�ڋ;��{�?o�i�q��2e�D�:�ݛ�*0�xӐ�|uX8�Q�9�Ғ���U"�b�؎��~*��m�����ey�)��V~�ė�����:B��HH�J���Yj����}3�B���u,ݏ/�����Mv|�m)HL� @g��7�>�,��0�M[�#��<�pj�Y��x���#���C%?�|�YJ�4�?�qx�Y��.���_�vaV�8��2ձ�Yq%��69a+��𣮭�+J���ȝ�z�J������~�$��{�p��Tn�n���rVY��}>N�\i����=�gV���2�����.�nK˕c��:q|0�8��$���AV{;�����0���@e�f�+%1���S�#��=Lٸ�*ֻ������5�4�{Gл���m�8P�e��ƅ!��?e��h�Ff�A&���x�c�a՚�AW�9J�h��AeZ�ؖ*&<%ua�t��CތS�S166��Ó,B^�Z�:�E-s�J���բ�Nf�>[�az�+���j8gHCyE�JT/OI�{F������
��U��VPn"�:�EW�D�$���+\x��]�v�3�3��7�.��Y�$)8Ɛ���v#����7���Nuȥ|�r��b4e�Pq?��Ƥt��q@��T�i�Ǖם��n�&,�>���E�J;O2��l$�Wk�`����s����%m�G������NLZ�T'9���c���t◤[�F�g���vPD�dLG]�Y�=�c�bX�v�U��j+a	�{[��*��,:�&c�t�g��$M,n[�uuM�����(�G�,��Q����˃m��@�~��W_�[�&��TQ�E���R�p*�w�&_�GDwWw�%�p��>dY'�Bg��)Y-����U+� ^�*KA���H����='V�ݒ��	6��<��<~b��]����vW��`ӎ�Or ��E�Nr��������v'�ql��5 �q �� �A`�e��
y5E*�'������D��MU�{��t�9;UM��@+HlS����p�bo�������c���v�:U�*�ꉚ���5���X��]�)��u<����oE@�B�� 
��}���J|���\��U�YR�R��Ü��))P�4?BH����b��܌~�q9�238��zې^�UL�R��5i"ag��ID#���1H�P�{O�����[A��~��a��J����2��PPiF6�5��QqQ��͌a��[Ф�J�y��P�]'�ED��S.���%L������3�_EB�ɼYc�L��������U�P���� ���yde��1\�A�=.�"ΓD�����6��]
; L�#�X�B��L/m(�\�U9䰦�<���Z��zt�5�+^�ED�MePUi9d'�X�HS?�	u�Z���ڣ�4X�W��ꬽi�^W���^b|͗,��j��9���)H,J�p��ϻl���;3�Jw<] {�2y_h�9��7��B�.q( ƜӴr�9DaB��6p�40�?ō�����#\�gt�ӏg�>��"��y�W|��Hi������K�}��Yۈ`-xMz/"> ��_".�}��0"��^�����K�<��͋@����u:��Ϥ9~V��NXC9UCf�&ؓ��ּ��X���>J��a0F�uT�� C�U`��e����w��5�ͣ��(��ϙ���,� kF��-:�䶼[�Z֘��_��ą��!�j:��Q;��-�mjB��G���FH���whT�i�"��p���Dz�����#3ƪQ;�\\�tTDK�y>�o�Y�D_���D��hFUU`_~+ڂ��FL^�N�3� a���W#�:,�. T����$��������򮼲M�3���{�	�|��d�[	��8X���6��y{��_,q�YH�0�. �AŢ�:���!��,'L2���t����lw̲�����S��s��bƎ��9��ɀ������+P-��f�{v���Ld��B�X� ����[���Y��A	o_9j�h��t`[,�݌'���-ǲ���ac4��%zo��`��s��L@?���q�	��(#1�wF���'D)yX Q1�O;�t�s�P�>�3�W��=my+�U�9��]Ƚ�Fv��y#�%Ͽ6����o���y��r6���ͣ���*9&�w�9�p���� L�ke�F�~�qPY�A�wψi�+.K�L�*�c���Ţ:8Et���2��1桻����U��o3@��J�1Ru��=��G�V5^�ؕ��,���t�|�N@�9I�x
U�~}s������t�k�}�ɼ�����ͯl� <h=X�b�F�8����5�l��>u���@	}�������s���F��� Ȭp���γ���2�- %�`���S�` S�c^�*��m�?B�ʌ��Ne�%�ލ��A�Vb-B'ұ_�Ί���APK��a�|n�Ф�SK�[>Z���H��]_9�sp���h M]�=fi`�i:K��$q���"��_�^�ۣ<l"`�G��]�+��$HK���O�a{�duzd[�H��;�(�S����g$e��?L_�ݫ��+g����<��{�t���k��tpcV�9xδ3�?n�#W�5���_�+u�����n�Uw�_R�7Nk�9óYJs�i$K��Q�tk �F�4�_1����iP�k�BC~.2���Y�[xȆLu�ܱ�j
�G>�:~��<��IѮ�|��=�[=���������4ǜY��P�T�)��"<�%Ð?w#������H��n2}kL!R����?��e$���M�@֟��ޅ� �V�",���b���޳u=Z�X�N�6�1{��̯X_�H%I� DS"B
4ƛUo˜�rV���Hf�7E�Qjs�/�.�e�o�&����m:�{T9�2��@��H�ՂUMf����n_Ry�혤Lnz��s�`�; ��Hf\�>`�N{��t}��鮝s��Q����r�������s��������`�\�|p��R�o�ג�D'B��e샄S趪���i6=��8Z��^��3�}^V��8A,�B�$�p�+�� ��?������p}Q'�o!Le�o� �\�i\��#i:����ΗWS��	;a6J�V�I�H�4^)
�o
��ÖUw�;z+Z���ux�Tל\���7
��$��8�Eޣv!�g|-&7B,)��"i��>p���ݠ#߉����_�գ���O��q%bUw�9�u@v-����+��`��$VǑ	%ߣ��6�QpPS�~�zE����`[��y)����!&�����o���$+lX�h��ģ}��&� ���=��z�쑾�›��˘swo62%�:���*eB�,R�P�d��`̠��?VWW������!_J^SSՒ��٠1�^�.��ʂPA��*�]t��x�53�KD���tϴ́T&�� ��b�٫����<�n�#؄N)�t��M�X�������p?!l@z��}���#7r�|�q�`u�8nK`�FX��&��]���M`���k�52E�Uy�0+��-�|7�:G��o�GhKХ
��BT��B�Z�݌y\��-�St���o�������9�L��p�4W�Rq�?*�ֱˌI���<���B��,��*���)��A�#^�U��o�7�����{�T�hω\<
s'��^kfZ���M�Ϋ#a�ό��1s�}�����;��N}�d}�%�zX%�&o<��ZX��E�Fe|ЋD����gu����"�Ӑ�Cr$�ꝗI��R�n�)�����;l��I��i��i��k��?��
�J �Q!fX�(��=8�D�r�
�;t���QQy-��<��	����6�f�F[�ļݦ�Du,Q����J�?P�x�ݩ �n�	D�:�6Q�h��?>ﶼ��tzTZ�����CB�|WUrm���_UP��,�aZf!̹�ջ�&ة	�g(��#��Kww�i�o;�����>1.�e�I!<H��m8�}��]�6�OQP�^D�Ҥ�����C#���hU�����>/w�d���Z��{������'�U�jѿ:�居�a��T�(�D<����(�v��:���NDO�th轹²�DeK�Y���\M��������@�V�L7�狾�2��F�=�O��|�=-�hD
��u�V�,F��@=� �:�-�U�P�D� �t�>v�K	è�	릊�lacm�[:�:��lf%���<ҵn������y�(��l���H��;�rWU�S�c�3=�ku���N������+�iON
Z�	P+��cV�ˬp�-⥟�L0$i[И s3��Q�Wp��pN��b����V�Rg�6�2%8j-���1a�fy���#v� A�^PCi>i��?H�%50O�a�Ѣm��ZZ�#I3��#]ΚQ8��C���y���4����)8�]|���K�z:!����d�����O@�;+m��k��3��-J�j�F�E^�_9���c�|6W�Sl��l�-	�Lfdn7�� e����D*T�{��~n�M`��{��9Jw*£�̑�'XE�~���o��Wo�]GН�U��O"�oMTCV���l�3뤦��l�V���(�c'Sʀu��Re��V�{b���ZȪ_��6!�V ��TuB�R�H�)�!9����+=�����g�9��c��I)��i��{���\�������[7[�e�e� ?3=�j)C5l�U2��$�2~�h�&y,vK�R����_Y'5Z\�Ƕ0.�x\����n��'{G�3��>��W#���h5�����4�>���)�h�_�sGb~�����Wй�rڴ�W�j��DM�n�!���Rol�Z�X�6~�� �0m�1w`�!*\3�
��㢄i��m$�7�hp��'�@�����y k�ŷkve�h����n���%SU��Y�:��r��Nv�K�U���s���<�������f5���	
��~=q5��VԾ���vd��<D�S4/�'Q��+�{�Aٳ-��	~�ۤnå+
2 ����>9�_����ƏCE�!V'ԥ֤]j\���GZn)����k�N��o��7�$�%�F�[��a,�W�[m�2���#^�"K�}��-���]�"�1�R!z���.��C%f0u��'���Čw�[B�;���P)�wX��� �涨G��C2��PW�fX�(�6����R�o8�	ⵒ�f0�D6� >���\hi�8�y�{hh��}�4���JD�ɥ`|k���o���[���j��rƂ��PW�I\�ɲ1ؖ���:5`{��m5|�K,���
d��	J��_�hឿds(d�Rя�O ���d���I�����ݙe�BC%7���h�y��b��s"�D�����a�f�M��\�_y�|:��<s�;�����3��m��[u_�,9I�9s_��d��J�q�a$>G��g��ޞ��>y9����|��B6�Λ?@���r|P�r�{52�Y�*�=J�>v���M}\���*�N�p�����N�J��X�_��� �F�q� .���F�Wjकl��nArf�Լ~�#�r
V���m|k���\Ǜ�f=��5����=���V�9I������3��#M���|u����o�I[
���1��m����l��6�����s��eD\�F�Ђ��9R� ���%��J���D�.s�:�{��͗��; �r���H�\pB�fQ$H-E����X��w�6b%{pM2`���:��3��9�A#�$��Ϊ�����['E��A&���ŷ��� ��QZGL���d6ɳ� 9޾`t1oCJ��A7Ώ��$$�TM.$v���p�W�X
�E� vp�+N�%j��\�`}�qJG n����<�����?��d��,�uD���F��뵅b��+˻fSJ��8y�mBS��敏���EC,�H)W�N$S�ߐ�5�l�;��e���`0NP����6~44�a�<�:_iX�w0mѰ`�4jA����潖�.��-���8˯8h$��O�$SP�e��ϗX�vZ��fkY~�v�����j�A��qXL�h̺���)}πH�)�����7z��n�7ت��zg�8�����07]�xh9/.+��G��FQ΋��>r\o���t?2s�)<�:�Y���d��.�YY�"v�w�j�C�~s!��($Uz�,Q��#J\՞�b��4�$���u]53)Etߘ-?6E��ߏx\>#�_2�}M�~�p�~(~�*���s��\�y?�))� ��ϳlg��wW75�R����4�дEU7k^sKjW���
�_�3���9%��<���=���z�zw 63ጲ�� �~�s�_M�>��1��x1���������@�\�W8-H�)��շ$�AYk�!>p�%��
&ڀ�30%b[ې�nە�t�̙l��L�P��u~��,ACǎsK	��t��I��]TdS����S����Ra$l�s �� ���G����)�d�YК��"q��?�?3���r׃��#�w����E��#�3����5��^� #-D��g� �����A�.6�]��&�`0:p1�L#R�@����� ����űnr�=�o)�a�>�I�s:Jr�]��1�dnQ��0���L�b���:x-��B'*l�_�w����E~@�B_�m��O�΋��@h� ���s��D
@,b�Ew�>4T~��EUd�JOc�e�OZ��&���[��{Ry4T�3x/^{���3k8�NW���]����${Fv\B��C��C���^᷑+y3�am-`r������2.F&7} S)�I?�~c%6'X�bW�bv��C�����P��Y����Aնm�r�j�8(�i��4�X���� �ӣt�=u-='g-�[ U�h�G,_��F������Wt2�ȍ�[P4$|<�>�w{���p�-fm��&�Bof1����`�6�J���[��Nu ^g���)gʛ�q�ɒvE�^�2>��h�qLV'O��vד���y���G�%a?H솥ӯ3`�"z�����[4��"�3�@LR5A��G.6��W��,k#�U��rz��wW^��76�C�zc����~�%<J� ��5�t��'D[[������R���)ߢ,E;3�4/�90�Sl#�b�ޢ7��|��ٟ���	�&=�:�T` �n�SC��Y��4ޙ��.:k��=�i�@�k�ǻ�d!p�d5C�^�J�=�F��[��c3�!7���]�,߈�=��B.���+7��jq��$M��+�n�{%� �y)��v��H�΃K<��k��`D��7�(�cS������E8š��Ю	4��~�`Ʈl��������"l��K*/	���n�]���sbrW��7#y�q$[�U��`������t�m�|�����v�4Y�v���������q�9�r,��Br9&��gTbG�E?��s�3��>y��"��`�"Ľ6��0i*����*%m+�����|�����yR��	�^�Q��josx>�°?Έh��AT��������h�,G��l!"��x�/�6e��/cvW�P8�΢�VwWb�e���$I�a���`��ݹy�Gf��(r�Tu-gHҔ�,�	*B������6V�@{��p�P����_�,��|�|���xζ~9���~q,z��t�3��Vq��;�K���=�y(��ܺa#������*�A[�M�#Ы|�ygw�Ӵ��HBQr���T�	���r�6����l�9�����[��%�$��W>j�ݴ�J�K��$PJ��,�����������q�ˤ�NK�@��ؽ���m��W��9
�m�~���*��²��a(2�l�󗢔����vX�5���ȓ2���>K��"V��$�1+��^^��X��=L"��c.��6;��*��tᎁ�X���K���$+SyM�m�H(��-N:���C�f�I�m�cq���W�zX�-�=�`��&u��|2(�Ԇa�_0x����̜ј�+�G�k�_�:��q�����*�xs��,L��ܩ<67�?�q���	=��z���F����CCm-�X�!u���Z�B$�F7�>���/ᄨ>�C3�I���ℇa ;;^�oMu}_e� ��ׇ��>�e�Mr}��Ә�T������ͽ���!�bR;ie�� ^�h�y��mc�s׫����M.A�6�҄v*����)!^Ga@�	������hiX���)X�� ɀ��{ug���!b��z�.?\^z
�E$�tFԟ{��^��5a�k�"<�jhDN�ﴐZ�h����$�IF�C�* �nD��E&\�^~{���2{��k��۶RDB�,�1r����-{�$� @qp�r|ώ
J��9M�����H�*vxa�NϚ}���<¶�w������E�mOŐ���t��
¬�!=g���z_n�ܗ�3�'☵����8�U���\/5V?Z,���To�zލ�5=q.F��'�9�n��Svcz�`�~��@��.��6\��N��V�3��z��U��#��<�E�Ům��Gq��N~�oOG�e*`2ӕ;ghd���������L�jC5P�Ȼx8����=�]�D���(�k�D�t7r����:�_�;=�@��]�C:2���.X�t!G��D��_G�"=��S?�����#�����ӻ��To#���:��|�P[�\��<�P:�^H1Gw�a����.��ǰ���B�qTR۷�g���@�KA/�e�_���]z6g��TE���{�'��C�]x�]N�ۮ���nޚ����9r�N�ċ������E9�i��G���v>�|��_�'И��V��[�� ��\�3�)m1�bF"�h\���k�'E�����u5?���4M�50*��K�F��by���s��^��(Ϧ�m�d��Ԑ����5Н
p���@U-�-�\ ��T�󾺬�Icv�w�E@?�to2�p�V�����������3@��$4x�u��>h�*���P���(+�N��㷄��c8W��g�8�U��8r��+/��Er!ϳ����Qe�L�!W¿]��1Q˳g�T��';]�W��K�l�q mL��0ʃt7�s:�߬�d__�V���h��#�#���@���2c���P1u -�R�<V�\sF����'���oʹ�7��;l(<�~)a ,k��A����$'e|
�b_�X�)8p�@�+T�K����֢��O��;|$۰��o5Xٽ�q��;�Z%�zW��Q�P)+u���/{g�	���g��NG��(:������:oX���,�hq�ˡ9ݣ�KtED�hV��?̽Vrr4!���ia�O��S��fH�����'Dsm.V��L�d|�n�ʨ�'���kK�F�ϟ�<V�Stǫ�V&�Z��^����P�ݸC��$HM��#��$����XT�)e:E!����,�t����8h�~���kM�	��a���OxA@څ�$f��Lw��������}��Ӡ�xl�_I)d1-U��E�;��5��J<��y�Q�tͰ/���أ먍w�сK�H�L�����G�Aa�����fh��Md.�4���eh�Y�쪳L���q��)�"�"��FX�Qx{�gL�.@-<T[���Ut����d魽��SC�@	�� �)��@C�	`/#�����P�fl�X���pJ�7��3�,]�����tXQHNN=��7�ܷ#��n9-M�-�X̝e�q1܇��զ~��P�|)B%"��K�~����N0�ކ/�A�@��;��P����Sk0�~�y�wS��?�֦V����žV4��&���$����.4,y�IP|�rl66�Q��7��\}m�d��*��V/ď�nD$P���D�垶�u��N ~0�Ry�p]YA�~Tx`�Z'*��7����I�+�V9�������o45!�A��I!�t�<�9'������r���^��RE��������_'O���PƏT�W���լ��'�g�����l] ��l�� �|��AA`kc���u!1�ů
�[)=DK�	XkI�y�q�NNR�u#-����V!q�{b��������5�������N4���_
|��ɰ&���\�&�����`��qQ��`�4g�o�Ķ�hY�
+�7�#sf�h֣�����)���~��C!��I
~	;�U�� 7ID݋'!��3����m�İ&TD��,�3 �ws���Ę��y���H���I$�Y=~�n%p4�/=�҃^�	ix�Dw�cA����1	�Ps�`������Ξ�5(7��LH..l�yN޲[�
=O��9��O�a�܏�������Ti�̚�gMH�$�J��>J���{�6��ᕳ�+�����初m�s����\r��&]-��z�&+0ć�ˀ���FX{�F��0��l���2G*r��4�9ev��#r��AZL��[&����I)����`�ڍ��ɥȞ�,w��}� ��9�ta�Iaڌ�?Lu�҃ �@|8ST�d67��`6���!�@y�\�y� d�W#U�򴸿գ\���Z���(e������r�6z���܋�W��_�6�J�|��ohCr���ޑ�B��$P�yK�[!�Һ'���=	��joc�5U���5ਣ�4�@�oA�H�S�ƍ�� cs.aIm:%񹭃Ln�1Ӌ)N�/k!Y��q� �;�K�л���C�t�pH�y�	��1ɎI��,��r�}��K;�����?�Z���`�k����&��h����D�{����ϰ3X�Ey"����}*�C�G7�>�+��5�{(���MR�<"�b�,\�B�A�� ������V9�{� !��x}��6�����}5��Q��X�Гp�\Q69��Ϩ���0'\xj�kф���M���e��D�����C� z@�˪ר�F���`2�G��=�B�x_�J�|}���zpu�W��B��w��M\�E@6��zS捋�!�P�
�GC�5���/3���́��j@�/ۑ�`�J��@��	(��Y�>_�s^�-\��DG��s�u�E�Eu .��SB���O�V��24U@����O��R������Ą�,Dѝ�i�!����A�]7�6'���� ��o	�RT�H�u ��;?���M�❡N���t����Q,��c���[�e9N��ľr:W��6B����\7��V9��Pg�W�}8�TT	+*�:�\�l����,Ӫ���0���p�m��أ���ᲆ�xʎ��5�V'��6�/����o��@_8ɕ1�K>wΔ匴����L��^2��cSl���/�-�e�����bl��P|3D����6hk?D�=I�H�fnpBϕM*P��H�h�)C��|o)'	��z��H&����&f���Z�r̐��1�nS�e��g>�t@��W��2�1����c�t�ݖ�0�ij��r�x�ԼƂ�$�F�?Nӈ����>�a(�G9j�e*@�e�z��]"��E��N1z�� Xr{4�?y�6 `w��&�[���OW�fՉ�*p�<X�M� ��>���ފ56�(C�p"IzTf��\��r�P�(9m�����ӈ�T#m0Wt�6e6�dJ)�R����5z�$&�e�]���AAz���&&q�כ9S�<���J��*�y��o�{������_�n(h]9�~
|b��4�R{�YʏP��M�G��ŗ��yc63�z���/(������hT.DR��S	t"ךc�$�����	O$���ķbѳ���3ێ#0��sZ��q }!��'�=.�c/��*Eq4xN/����i�6��6�#Sz���-�MJ���$�_��\�,���tȲz����%oKe'�ت)!w��}�=���询�:~M"��&�;��|��w���?�0�vC"����WĲЀ�J�#S�������"Υl�d	y�zh��ֹ����Ըp����s�Fy��ḽ��3{v_�Gn�e�r����8�δ~�XWӒ�Xc78*\����q�c�)j�L�O��	��e�E���
w[�n�&]L�>�Nf��� ��9����(%L񨔙�;��=�d�*��_^�!Ä6O���ܟX�P�6����"��8)J�����U�3��f@�C2x�P^yn���g�����e�[��\�]U�[.�·eq�Y���<Y�Y��d(��ɰr6ơO����r-�O=�$3��ǩ<��lvJ�R���ݗ20��S�?��>������������z?�̾�h��\_m喲��ԗKa��5�E��3iw�5��V}½�]h�n ��𯛼�y|���7/���@�A>��Z˭;1�{��#6�tox�O�r��2��� ����#z$���R�F������	J��A2.�m��h;-�Q�ig��<��F���`��~E��� z"��s}$�ۏ���Hy�_%��'&u?�"����'����6�%�ܓ2���W�,g��^JO��E�V�cj�';��2��ݑ=?幃��tY���r.i�"��Ýx�܅i~�I�-@}�@U0�ʌ�9<8`�HDжp�:�~��]ѳ��I:�i��̨V]�d&���7�w<��ӛ�� �ϓ��9E���2�X>�� �o)ҿ*�DРZ�W�[k��=��#�?���~�"0�3	p6�A��v7Z��d��~I�j�
E#_���1�d��ʭ�H�%7��z��9q�.�m�I�o8��zJ�xϨ9ąu�ė���˶X:��(��~ξ����O��Ϭ�&��G���T�-� ��(4�Բ�@�L/X�o�����r�9V�t�z�>8P���Ķvo�Bh4@{����]M\�+i~�"Д�0P*�S���B��1�s,e�ߝ㶜�aٗ0r�����?���[/�ɋ �3J��8D�t��m���ȝx8���U.�F_w.�]���q:>��%�iI!Mggd?K���*NO�����m����'}��f�sM�' �b�[o���IaE���T���h�E*��	#��R����0i���W1q~��l:��M��*�����Ի���4�w!� ��絋Ȯ����>	w>%�eGǗ�2��ް�B��I	�*�JT>,\?�����KA�c�y�P�/x�Z�� ��/��J��Y}��^�?g�BX�Ə,� ɫ�*�I�o�COk����˷w�w7�! ��˜����1Dȍ+���6�{w�s���+�T�-�^�\�x�nR���Q��e���|�Ů��V�[2$S����%���[���1;U��.�?-�w���-�L���{��	���/<����TtF��'�ڔ��E� ��f�Z����� �ܢt"�Í>��h�?'�5�('��4���f���xoX���f�i���P;1���`�_����-ȣ�G����BoKY���}o��Ɔ�	q����*
���G��0�~����ʛ��-����T9�{Iнw��sgS�ixPf.ݳ(��K-*6X�_�bs�����1KO�)��@�ø͙��*װDc�H ;H��A�� �= �?�I��z�{��:J�YƲU?�{0�+4�����C-�[��i��ƣ�:���2�Y��o^����W/jhu���Wx ��ʆ���,)--?x� ���<ڋeG3�ɯgm��A�ѱ���%�:]2J��
���E訅�iF�J$e�5�-=U��<C`�U��#���NR���5.�.Ì�,ռ3���$S�G@C�养��m�dz�,��O����D���?�v��N͊k�duH[�f�8g�"��B@��G�������wj i�r���;@��L����5m���bLXeL@���C�B�K�s�b���l:T�(m�A���;#�v��PabۇP�<�К*������z�@�>�t"�l��P�E��MߪR�z��G*�Q��%�a#�f��eO���������&d�eZ���_ 3�q!�8SZ�[Z��k��\�c��0�u�i���DP[]1S��|��ٹ�	�i�v���hȲ/�L��G�0r�8N�93���	��y\�G�TH���c[��&,�f�R$�
__���v-4��E6��mъG�P|�<��so&��=?���T����������k�a~1�6ɛ�G���b�\���!�B&W�1/� �W9U��.��h�����4
�(>�N�Z��1k!:�X����\���+��l��m�ܤ�[�;�9ѧ��&��A;[��b+��7 ׶��>����p�j%�Pc�K� ձ`G/�-��6�`4X�yw��D���B��N=!'�c ��p�J���߀�T�w����2y��;ږ��Sn=�8�%6V�7L�J���)VO\�Y��n�Pb�fJ݋ˀ��V�x�Bl�����1�9���[�{}���Sği�q7�Z�6���֡�Z*Z�c���%~���-�_W>� V���f��P\��|��
	��04ę&�:#�e�'��B�i��SY��@�0��n��=�Yإ%_�F0�(�g3P*w����O��Op�pѦx���(JhT���D�e�k�+$��G���1��e�Ja�J�I�@����[�h�@�R>2�,��U��^��<%�����g�/�hfe�y�a�g&e|8�2�f�[Qo���8��
�0��y��f��>2_E���Ԭ�{Q�k�S#�!>ӭ�;MOn��ϣ��j�ĸ��2۱���ɀ�c���:@f���zB���J�:�g�vC]K��=T"�Y�a;"���E��,u�ds&86Wz{�[}sGT��Q��:�غq�����;-�N������~��b GS�Y�:�N����<������w4-��8��HG��|v2=`�bՇ�v��)v&�}��:��@0�.$R�y?�x���so�w��V*���T��/u@��s#SXI�����IPz���Ù +s�(�o�%������t��C}_�C)�p+�����f�i�q�����S����ɥ�����V053��1Ѵ���y��$�V�H@�?��7����6Ͽ�sf-��@�����A��(ms@"�s��;
]0�GS�;����I������a�y�@vY[	�U�6~i�taLW3O��������@T�~�c_d�%:�g�V�S�yRU�2��<щ�����HԿ��F�ф�y&̕g���#QBܔ����$���)Wv{���M��F��,EyYz�"�
6�$P)���`-�@鿌��M>M�f�Ow���)�\�s�P"�β�"�����Rm �u��I��g�E���Z����
8h1($"�([1��(5���+��� �ri*rVx��ȓ%N6�IcY���b�_Qf�{i�؀E5W���S	�U!��� (P���J���7m��[�Xd���Q��#�s�g�� ��к��b$�3��"���`�4����[x�/�.L���6����i&w@J>>uҝсz����Π.H/X�r*��J�D�#?�w�o̒_�V���@V@����xǨ�S�G;�U�9����{�j����>~r�r�`�a��ڭ�� \��g&lIu�_�}�9JJɿ�wC�4�aυ���H,���'��90��7�rq4bH��t����aXES�I���@�7�U�dLei�
7��ds���h0Ϯ�?�Oc�iu����r �K_�bj���KhL��!nD�����,�㸃z�|�ʌ��?|z@0^���B��0g�>\�qq��5v�����kB����Co��m�:��Ti*����Ő�y�$Ea=��xg�2�o�G�I�w�*-KwʭLf�թ�ՠܷ�x��;i�}S�����+j��u�S�R���dp٧Y'���O��h'�G�9J�\��{�8�®TJ�c�)����]�Ѵ�9e�-`v����� �ou�`���
.�OZ `���{X�D���Q�a�=h�̼������5o*9��"���sP/�I���@��H�y٬l���Z��/���.�o%�����K��j F� )�Wt��*��=?�b?B4Q�_"��9Wｲ�������� -n������!fi*�����;�)�	6M�C(x��]�+�3X���˫.����bӠpm��8mN��f�ƥ��A(�o�T�(7�[4�;b���[��!��g�!�ī�VZ�3�h[�k&)�$��>~�=�W(r�Y�(0��}<���p-񏇗^�_̃CQf�'��m'��[I�Am3����gq��ⴿC; �����Ȉ�+����^���KH:��9��ν�����&}�X�I<��I��J��t������x:��R���$�'6�նD��0iQ���y"=��{�HV�'�N���߀��a�`:��i}�紛s��N	w�r-�̰�,f	��W _��b��u�E�ʕ�.Ktl�'�3�$���ƨ�܏W���%?�E����k�U;@H<����y)@��7�&�W��<-�N}���^�Ct��(�8��"uV`ѓ�(�_�H�ġ�w.��U�d�U��������,C?�5���G��M����l�S�1�A�f��f���?+�9��	����4)%�Ow�ސ0�=�ţ�0g�{�C-i�P ]����^���&W脽�g/gW3=+G|<�N�6�� {Dv�$�4a+�H��c����$ lJO���ڊ7% �;ٴx����rf�?�?�jקs>�g7��֫:���H�EX�����l��9 �Fӽt��y�����*��> �}�I��fF�	��ɳ#C,	�xvus$Y*���?�C9���fy|��(�6�N�)���oH�2x���17U) E�(�wH�y�\^��٭[͜�O�gD\�����ʼp9X��7�o��[��P"U<�,|���e:���}�x{F���Zg���aZ���}Б�y��_I�!:������]����\�3�0�t6 ���ޣ'����(�97��k�������0,�d���xl�0�=���;V���aS�&�,G����M�Y�eӵ>@&Pą�:�|������]�v6[�v���y���-�U�x����;�Y(l���u>�m}�;��U�[�;���)��)��\"��Fc7�`��fO�z��pj�Tމ��$}}��sK������w�,�o�������귬�51*� ���	|g�X�Jd"Fq��' I�\���
�F�󰓠A��'�E(�h��2���|E��� � ����Yk2GP�e��(`��|���a/�X��n��ʼ>`��w����u�2`,��F�v����7�d"����w	��br��iBh�跻��+��j6=뛾���9�¦�~�v7��N��.(`m�f�R-��D 2�9o�Eg���7�A��Z~szc͇��+NS������������pJ���~<!��t�(�\'�lf܈1�@��7:�5���n���H�=�'�
sk�����e+͕��P�A�F��i3���q$�����*��E�e�k���l�6�:����VI�*H�B����
�S����x�UrH����~��TK:T��r��$4���� ��
�U��xnZ~XD
��}�y���.m^y���Qc�_ݴr�-�4�YQ�����x>L��M��r&��� lЬ|�x@w�k.e��
��`)�Ȝk.l�h�eUd��\�rz��X�=�2x�,�c[�<3)��C`�:!�W\�b?tj�~�}8qt�Q��ɞw[`�K�;J�H1�?��^q?�rV�L��V� Y�����K���dii�V��f�r?���*���.fv��O.X�\�w	�*j�Z����w�^p��.*$�j��|�}��)Mvk��f� �.�����X����ֹ������R�/}��r�P�ҫ��LV�~��Sk���D��4S�2~\Q>��HSԄ,�@�g��3*��v�ݮ����D��gm��h~:�V�5n?�4�P.cn������SZ�y�;���K�Z���)�O�E���u�Opتd���#Hq�wWI}��j����* C�W6��0�c���} X��)d���A�+Q�o
�}��
�o���j��n+wN
�q�;!|�8���b*���ü��ٞx����f�u��k+z3fq�{h�2q��x{gS�O:6-���{�?/���O=����$�;!�#(l����B�&b�����44���|�>��6��Hr�Y�X�js/�!� cw$f.k۸�n�����G�t�z)���x�8�Il��Q���\"�� Z��E��y]�G@���
"����
��ٜ��u�����k�cN$t�<m���#����
��bҜ"?׀OkyCyv������Y������66s+�{YvaK|�&9�� �o�l�O7�u�q��H���)<جp��*0o@��!o��"��A���fX�ƀy�xI��"�?�9�c)�/���۔�q/�F 3$1�\�(�{.
�_e�np�E��{�O����0�����5hO=sk�v����6��k��vM� ɓ��Z�,��A?�G��M?/�8�;4lˌʌ9��f�^�FL��r۝�� 3�eh�t����.<~�J4���קj���Ʈ����r�Q�`..<�٥t{��s^�����(r������WV��jg�>;�Y��S"�6�H!h}����g�+el����E@� �f���"2���q�EI��1)�Ԥ��Db�F_���VA�������Z�c�n�U�ҏ��An��"�ƶ���5�����zt}�aO�2H����Xz��a�H5��y�W�_[Xo6�n����/69#aT�f�*�Z��*�k�0�*����)�v�sֵs=�=J��p��w�Q!e"Xn�r�E{c�b�
&Z{�����Χ����ɀ�k߬�v `�""��
Cbĝ�S�f�U ��[��J���\�V��_~7�5���0�Cf��KQ��4��p����� wb�M���Ī@C"�a���>���La���owb��"�{�m���%u�c$-�j{6b���q�"j�_�.�h<�W��%�	�Lt��q�uac�������b��r��hS�l=������c�Z"��5@��{)n��1����[�W����z� C��&H\\�Ot�2���n[���l}���w�_J$��
z�d_�YZ	(�kN���JXg�W?�_\�W+��oЮ3�*�A�a�Z`�u��~���\I{L��JMя㜂��C:V̍/��ȩmvx��vy��rE?�H�sݥ����}H���E�rT뙖>>l(��0Mr����^�g <S�!gbB��i�������L.�,%s$!���XEA
B� ��Q�<@��w ��Űdڸ�봬*|���	`�B{u�L8썟������߄'��y��6��� ���x��/l>�3���/�GF��o_�2����8楍J��k�.HQŐL~e>����|F��L,9��<�!��!P
�5l�c�p.3��r���c�
;Zv��\.�3�n�*�jR��v��v	��+BJ�+�T�զsk8������:l+P���RK�;��4�����KFU�=a5�(��@� �*o�_�Z��������_�xz�{r�U����t���=$���&W,\�fy��H 1_d|t;̐_���t�~r.������xHQ��E�s�x)�h	���++��6g^�w���X���hh����m@a���"O�hl��PO��X�x��	pvq�A�ӝ�T�iS�6&Tʍ(7]~6��ƽw�P����t�<�BQ/��e&���i9��� 6^�$2�u�,���m%��՟�V��ٯ3�c��E�N-(�l�:���-�1�o����@q �톷�b�e�zA�d��T�����s�f)k_\��k-.j
=T��i�I����-��� l���W���{ڗ���c�xp������n�0�p���(�h^0Ùέ�p��a��j���ЮP1�`�蛕*����r) �x/a�k0�}���BH���QIy~Z,Ѫ��P:��1!��1�9�K��ݎrbCڌ�h%����ѻ�����$��"��oF$nꦛ��<���k��"W !U��B>�Uд�j��Dkʬ>Cr�|�ڧ�cm�� ��{/�Le5��r@G#�|ܽ��g�9�*��o�n��������yN�`��y�t^�}�o�S���emLJ�����K�Wx2� ���}:Mg�U4=S0�fG�ɮ&(q�b@��Za�38���!��w���ʠG��A ����@�R�6F��t ��JAi�W߮�A| �IM��6� .��o)�|�@���a��@TR��Mٕ��|gE�3`*�1|�/o xj�l6�P�?曦ĳ��	��mN�P�<rL����\��X�W��Ts�HDR�`!G���Oݱ���l�Y���_waw~�;���a+d�R�x��4���Z8�ǹk�]�o����q=�߯ΤIc�����W��UR'�b�=\��O�I�/�(bg-�y���`lwב^�Ĺ9���*.�LQ��{U���yq¹��'�b(���;�eǏßdu�������_�}�?�����:��ڷİz�\0��*5�V�����~�3���d��5v-�l4?��0����j�S��N��-pйwN�7�ᷘ)&���Xӝo`ɂ7S+���V�Z�Nv�m���#�@���4
�
4 9�΍�(& )�'�����
Dud ��w��ap�8@�d��S���7�mԻ-s'3�YN�2T����N�34$�4R�ʒ�Ci�jy���Z%Ӎf<	~�1���:,߭�oc�Y�	�����(�]A��g��**�`��˂S�r�̴XDЕ���p��P�y6���d|�fݗ���|A�����ՁA,�܂b��!N��з/���2�����Cu�'� �Il�B�K�G��/?9))�-a->�JBW�M��+4�n������_��i�Z�����M#��(a�L�#ड़8�R茣#�3�0|^ѩLxxy�v�7���QÆ 4������t6���QS�l��&�_n�F��ƪ�!$5�`�A՝�;R�dQ�)��LB$Mx��#�&K���<�Q��`Ix^�C��N���Z� \\����	�8XY�|ժ�_��Mq#�J��>��]E1�-��T�<^J9�S;�r���/~I�c�ܒSj}��wk�rhuȉ���Bbʖ;�A�b�ӛ�!y�Vn6j�%-;�� t�h`��?>���p���o�Tp�`�y9&K��/�E��%��_���!$�\�:�\���3mWa���N�Q�_fd�C>1���jJ���b3?T@/��=����So�@'��:��lɛ�9��B2s�ķ�Z�e{"��~!��Y�u����I�T0��h0P�)n?�a�v�O`��aoM[5s�J���}_17fɤ׫'a�C�����d�^�x�G�c \Q>~�&��?$�z/~�`��]����j�K�]eI'�I�ud����I5�D%�r��ć��@S�������m������y��۹a�+?k/�lm-�?��C8�o����w�=�IW�*֞�d��kP��Z0��n(�[<�x�P���о��=�s��M�U��f3���+zw�������
e,�G�a�b.q�[���NT�#'�d��w+ ?�jnc�D�_$�t{^%5~7>1��]�qc4���uV��G��LV�-wB��2v_G����4�Q"�/�bX��5���S�]S6��罊~3��1P2
D�!�/`'�%r���m0xɜ�HD����w�U���!���rRd�$���H�[#����S)ڕ_�XgP:愑��Օ�拾m�^0���r��^�R"�#{�ܮ�e`�b`��Ye�Z���Ӯ�� ;��0?j�"	�ͣ;��D�9�Hv�(XS�j�hw�D�[ *�o���{F=������.�zM6������1�����g���ڭ́H��}�=�#$���EyoV����_�u����B��*�v�{�	�P�"��)�~��+���֫��܇Ho��Z���hE#��_�3i�%�� {����Z�"D��0;�o�+�$�1w�y�Q�y
�T���J��ָ@$�q�n�z3~�/{��I�5[t���'e�?�Lz(aO@�n�Ia@���
��#�˭ٍg�	���~��?������sז��d
N�p�7O��m��~+aV�=w���t�H�1�����4K�����mxN�uW9�7�L[rw�OPןA���w��L���gS��&�IRJ�z��QL�U#nC��Z�\�e��d~㓡�[��?fv�߸0\øɮ���ו\�i�k�5rqkk?O�3L����y�><+Uċ���yӘ���f�6����L�`����xqaѠX?���:���!w�R�6�f����.�Y�ދJK�l�u����5X���"�x���wOde���������d5j��B
�}�"/�'�{�+>��n��(�λ�|��wt��4�«
�A,��E!:��X��(�z����*�t��7�~d��Q�d���8���J�~�	�!�ӏ[��=�|�2b����KJ�z`΁����$�iC]9�#0vpD���£T�����C�>�3"9*�4	�n�����F��JHe�9�z~=1cd���z+��3��M�6�CF�ߏY�-w�D�#6��؏�
>>&@9���yy��6�
M�W��M��r6J'-�8�O��^��;(����r�sh%!%����[���ȰЍ�f����7^��cړX�޽޷��m���~V9��E����c毂�棗�'�_��:'_�*ݥgM�>��r�<N�>EA 3����1>NK*E�A�	�!�o�35�4/x��U��L�*��E��1�؂-`�+C��8?�R���ܞ~/t�k�p��=]J��q�F�����RD���� ��� �W�PdѨX��U^���r4���k���-�����V�_��|�=�U����:����~��I�)�!��k�_��;4����^�ƭr���W��N�&�N����OQ�+�F}��*|�5��x��>`'���W� ���p
{��D���UzCX&=����T��D�@�HJr]�$��_���jإFM`x]&��46+�\{`�[�3r�4BHfl��͊��_\8����)іWϺ~$K
R�!�<IÔ���hfC}��O�-�T�6��{������,�(��ϛ)3�r6�%d�d��40OspЉ f����� �N\�د6�����G��@�V����*�S�ٵu�l;m�n)c�;U�7r��׾'��I���N f�����4�u��R��V��uL�ƕ��1$H�R��.FN�n���-��%�QWDF��� k�*�Vs���vKu��H-	�ȕ�� t�Sm)I�C��F���I%9���ewD�B'��a����ž�z�I�y�����y����z���P��e�.�a�~\���W�]���#�5\4��T4�r�r��Gc����O��x���⚽�攂�\y;L�!���4#�ۿ���00�3p�"]�i�`����]wn��g���8��]�F�! �}�&������-�r\k1�y�z�HZ��o=h;9��Z�Rp�C߫\|�*���!��jN�'��/i_+"�}�Z1�1�&�Î�Ï8*L����wB����U���?"NE�*����28��M���_Z}�A�V���>���V�5���:�C'�� ��Qt�(<�:�ԾxJф�	B
��NY�x�9h��s�k�4"���V�d@p!?�1F�I���\cˉ�厧_t����t�����w?��A�?�O��a�9*�̒�XP���f|?OG����c��kߔp����t�����Y,ͮ�1���\o�� �d;C��]G��I�lC�����v�R6�7MhSf�h��RN��>k �K�����2ǌ�����"�Ө�ٽ��^X�Hr�|��!�kM�x�q���Vf*�������
�}G�i@c֤���p@Nڹm�������
T�&�AeB�P/���i���?p(7�z��0\^�;��F�y�ۺ :b�%T�M�U竐�`����ն<�^�*�*c;��T���nٯ�Z�M��'Ei���:�ӟ$�v8 ��6��بx�K�BX�j�����r�.�ws�� ~�`r��ᤗ����js��ɤ��X\��a���ˣ=}VV](��宜�<Eȷ�AӲ	���4	.��|���T��+�,0�w�bԣ(�k����@�Z2w�(�z`���T���e�(��7�0_D�/���*��/{��Qâh��ȣOu��99��>"���Ճg���Ihƺ�qp�CK��Iu�ٽ����?��)'I�@AN/=���˩b��@a)P�ˍ��4�
�F��x��,�P��8�}$�� VpuU归κ�}��\�>�Oy�Hq�#��#�5;p���SA��w�&{��`��=��{r=h�\��or����zmF���7�Z"��%iRF���^��K��
J0�s�b��m[������P�*��To�Jx��G�-4e�-�-#��vI�"$���
_��g��vǑ�7k�j��rS��5,H�2�	�.�0{w��XVuޝ-y^�8�e�� ?������\�YX
*�N�8�2W��1�Gʈ"��e/s1��\A�Ż8I��)5f𦋿�a���m	��pYoIo�'��4Yh'É���\������EwJ���2"Zw-�	�?u�.?�[2o�t���o;���8 "�~�ߙ�)-�AM��R>�;�p=�cV�j+����`��4��m�Q�@E��CCb�SI�P�i�T�GY������;+I���9m�T��|M�EQ����D�7�3���)�wT9Rw�P9`̶r`P=�9�@��2���;ک�\�iwx�;/dG���^qFj������/ń�g%���=��c����1�`Y��B�����ܲM�$���mL�߷ն��{�;A7!���������Րa��u���67��Ћ�dZ�oVU�=1����o�W��C��{d��3�6n<����f1��1������G+���l>����@�$5���7:�!��@�k�k�e�$��� y�X��fE�Wڛkk&���k>BX�`�&��c�{)��rz��R$�B�r��fk�'��=�J�����/蔨d��$�4��3Om
x�H��qWA�@��E2�`?wO��]���n{`��x2�?���\�>�o���t��=-�ǎ��&�\y�4�i��[�v	&���κ�x�����+�4�s���x��!�����t�Q�h�} ͮ�����z}�`�1�p� BQt�QKBCw1w�7N�F��D)e>���*�Y�̱��/Y�q�t{������4/��M���D�z�/������F����;]�Q)�u�Űƹ�ӛ�;�׬ ��}�-:�
���<�5�!���
-�C���rt�>ê�*����c�}:_�"zE��U���)دc�>���p�J����	�;�Bj�B��;��A{?'��S�徴�1Ԅ��^����nz���(��j��!�¯�*�Eh�c��?.�=�\�h'F`l�THJ�z��pR��v��ڴ,��Is`.�o~`Ӡ�Ky��ǃ�bq�����>I��˾%�&5�W��?��s�������)���O���i�����x'@���+�c��@����~'�$�v����0o�l|�w�hQ�Y���t�+� ��!I����M?�{&K�8��a:[������Ȟ��9�QO��UI;�;Ti�jR<�	w�OTJ!W�
�;ō�����X��_�Ȼj`����P����tog>fu@#k����H>Z�(S	��"�@ �$<�Kk�y�ZT�4�b��VE\�w��%0r���[�%�F�x���D鿝�b��?���n���
1h�fڣ;g���u�)��cc��md� ĤN:��n~�BM%�8@b��������Q|o��;�:��Rr(4���p�ԕ90)0�E�n⟼K��O�՚��uR]��j��/�7���)�?Z]��J��;��$T�2�]ᣖ[��$;C�]#�|2������g5���
��%�!��C��&�t�X�a߈5ݶ�(�iJ7 �(:�@�Ժ���c�
����c���Ͱ)�V��f;�%����Q�F��=H��ĝx����RU�NM�޳2^��ܪ����ȴ/EYg6}��L5#���$}sd���G�Sj�HA�����ٿL�ִ]��W�0s�J��)�q�((ML+�GBq��ȌI��2�x��Y�С�Dl�<��)�Q�72̝�L\�v�ԛf�H��,b�[�N}��dO��e��ߍm��<��hd��>#.i� �E������(~�*�#?xQ�"���Nb�x�6�Y����:r�q��`<�@#*n���խ�p�x��l��y�dP�Z��9@�g(� [����۲�ͰE���lJ��c�m���8;5�-��ja����Oo"���lRp܌٘;n���*?�j�|j�`~b�2��re��D�m�نW])�lڳ?�.$����u��~q-R�� �c�y�⫫�J�#�D�w�rc$�v�>��+���W�A�_]ܱ�����*\� ^�+�����['"���+FVH��X���Q��4���Ի뫝��j�j��z.\�d�ӟ�����:����Y�3��JC�����E�M�W���j4c��ejixG�^J�)s�ׄ�k�X�S�8((U�� (�^��s+Д�� r��	��� ��&�Ĭ9�g�'�L:��<��y+f�����¡S]��%�j�u�hj��E}�,`R��d�k��`){߯��H�ɠRC��9{s6��g�}
�̴�#�V����q�z�A`�$(Pڵa��/$3@>��|��K�|L�tw8|PQq1:���vn���W����o���m.c��љ$�ò~'�΃,$^��ِ�#guU�[C���b�1�⟎C����L�3@lڅ:�*Ye%c|�n5�y�<�6t	?U
E�iO,�;���pY(۝7��f�¦k�I߼Ҭ�}oKf%B�r�w�x�$���nx�S��ƽ��#�]�)|�al1t@|����Fr���q�aJ��zT�k����|p��2��M�5�~kD'���8��j�hiV�`&o���K���94��	Nѣ .Ω���3vB�aFJi��OP^��;V{��z��u)L����9�;���;��J[����+��p�.�Fiәm$9��䷻��4ɧ�����;����F��ʘqAI-6�V��A���m���\�=�s�
^A8�nz��~�/m�a1���ª�}-�[AY7����f�>�_�d�q�����>1�L��2�Fq�Z�1_#��Gq}���Ћ�2���4Ly{N/&{w��N�Y���		�"�i0kjY#�[����|�;F�.߂i�zh ��9�+�0���Oꋏ�[V�����zE�Q�Gp@DW��U�O��8�;� MM���\�� H�[(�t�y3��/lX����C�-���Ȁ]+t[s��YZ�5ҋ��R%��
�L��&&�p�n{#��]�C�(���2kt��	�/ϐA[��ؕ�:�C9���a��#��K�u$$��Z?��e��Ԙ���� CZ����pK$�x��t�F�jiP��M@�����&�l�^Q.OU
2=�x=�M��^�:����D�d�6ף��sD�2�S�W�0 v�}��J����M�[}�/c��IF�����(��!�&B{�v�R�h�	���74/�h7fEL+���vP�V'��	2�}DB���L����i�JJO�N�*��$ɤGȝ,�r�$|&���X���uU�~G|�g�^��0lG>uY"(��>�!��\&�@���(X$%��X�T��{����4�ͮ�C�	S.B�HV�~d�$���8]f?%,�s0*�Qe�/X��V�P�`g:����y��մ�<NF|[߆���x�o��khI��LI�v�lT�S|?0b�"���H��iv�$wB� S4�fO��2b���y���=�*�q��̤=���0�ؘPW�`�OT�w�����$2���R�4��#�:���e-���0>#�MZi~����c��1[�P�� V姮0�WX�{�|m���ʓ&�a��U1Ξ+�ٍ]@�����
Z��!@��}!9�`�|Z~sNMUa�玎�����\��>��&��ީ�,��T����q�f/k"ô���Y�/�Lљ�� �Ov2�=�ən�SH�0L*-fz3R�&T�94O�z� ���-lg�1uڧ�v���[�m}����n4q-q[{⽹��tUC�p�F�:]ڳ���6���\�*�v���G8:`�ȁ���
�����܊���wto=�5w���;y5���/q�������k�?̻Y>|Pl]�H9U[��5
̎��;%5=�y}���4c�6i^��O���DZ�a+�mH�ͱ�6	JXl�j�u�r͔�y���<N����;�jDy�iy�:�T��&tE�	�vT<b��]�n�ꩂ��=��5��c�J� ���D�^�Уj7���}��Ӫot�SX*^uq����ıe����us���X�-f��
b�/้5�!��{���d�a��h�X�5A}�vK�;��x�Ĉ7�����[�y 4�=��v�g	cQ�N��Q�DD�M6����(=���7w�\�{4���a K� �)ah��j�tg���3*�nhe�v۬9��� ��a'��p���YB��Ї�35go�X�������f�C�WC�K�U�6�o.��u��Y8I��!g�!��A��
m�>��FaܧUWsگ��j��4�;Sk�2`8�����o(4��E�-ZS���`J�R��b����K���E95!=ߴ��t���i� ��T��H��u%R]~�ގO�ҝ�$�� ׽��q�o�[əR���(踙��q� -?���j7.^엙ٹ��whf-�3��P����g*a!�Z[�Lh����X(��yT��o�$3$�G��8%�A냰��J����$_� 48�s��<��>�$&�k͡����idQr�/��H�V���Db^x���[� �Ol#r.쮐�����]��7\gӵ��x�X��kU	cm����W1r-9�ՠ�#�h�}�ǝq��m��F����̓$��$���G����5�:�ي,�YB�; j���*�� T�pN���S(<�ŪҒ��Us��;,+g��̵\�
��0������of܎��Δ�ϋ�����X��2�g4q�.��~EAo{�3
�m��so/��,�'�+�x�<�;?�SUb{�QLО�g��`O	��Sˁ�K�{䰯�+c��ٍEFYjG����T�ɡ�_�C"4t����FDO�x<o7���$��ح�0��Xh7 t'��/��iUd0�~ay�i3ͅ��'
�C: �K����&^ʧ�e1N�a�v��c)��Ѻ���7����;��B"g$�N����&�~&~ʤ.���|J!y/�C�uDjr��6�v��k������[H}+��B��r���3��BF�{�k���Ԛa1�SY_�Yq�B�%	��oKzD��-��Q� �B'���'�Q�Y>����=�M���c^���)�A��������	�dsd�ݫ��
~�3�NT���k=��5�mx��5�
�4��,9z`=��{MS%ͦ��/i�1�_ C�Bǂ���2$�^3�ʵ~�.���0�WXm��?��Qd��0���,��CDl"""]z߰\�Z+��g�͕��& y�n�[�v̘	}5����F~�s� q�x$�y�A~��V���
���6i�g�u2���]ж�xaAi�+7�ʨ���
�)G�U�{ň�"s�ׇ���W���.Z��p�6	c}cQ�>��u�U@�{�WR�P�/�3��4?�"��� ��-��C���=|�
%ö88��r�!b�b
�{#sӦ�g��������R��K�<�L�u_�-�a��"9{�:�*N�ZD��4v1 jM��W��ަ#>�`�
0z>��K�v�.j��E7�m�eĀSk���9��du�Xve�4������I�w��ʃB�O�ly%����q��. ��� Ė�������x�#-�bE+-�o���|)C���߸/讏{�ּh���h�0�R��
����v����D�P�E�,"ZX�AN��b�����'�)�@����N�Y=&g���Yz�gV����Um����)���L,O�)w�7^���}�׼��� 	(wF�qn������& ��T8�&3���u�`��2_"����|$���r�|�/;1�����D������o�<_J�k���.*�V&ba,���+�޳\t�U �	�ie���V�H�����U�-���S���(���
`�,�ٮ�	���9&�ގ���֧��=��' �l��N���p;!�������]�t���Ȇa2�Ϊ�}wG���|��r���w6�����(���l�x_Hg�c[�c��/S�W�JD�`�U�{|:;��;:����y�ڈ���Q#=���8
�r7	�O.��d��3���|UN�X?Pe^�m��qf̃c���-n�X�A��~d���{�.�� \��G�-f��v2��;@m4�W���.�.�f�b�#JZ'�Kiv�\��� �h1�1U��&�S7�'f�~��gR_>:F�;2����a�n����g���}����nT�Q�j�>]�U�(���:�ؐ��f�i���$��)>����DM���d�������GW�����R*�����WL4�^u;�cv2ABt�ҏ�*I���~��/8",%w!7��J5^�4���x�����\��- 7���X6rY��N1z.@�%�=��5�N:6��I���0��9;� RI\�2� ]�`�|W@�X��t#2���B�V���N�N;*^��q��t6e��>~��F����"�x=���?t�ndW��f��^͇���K��i<�xl� -'����H����Р���Gp�����7G�bn�1�ۇ��]xY����V�(��JѼu��'L��A[5}m8��l0f�~<��D��!K;��aꕫ�� �wt��y��9}d����},��q�qї��Ɖ���(�:��<E>�\PX����ۺ��ܙ�Gn��}U��'oq�7!,'pH�pϙ�$y���&MB��������Vk�1��B[���/�h�C���]�Kt<�$g�W;=k��1�M��Kv�W��+��'�L?����H���1^J�lb�3ꪆU�^����*���, f�]�nC�6�=��C�
��!�񭪫�->��Ĳx��[j�AT>3L�2B�~�Ri��q
�V�`F�y�!y�0Da�	�ڿ����RZ\a�_��S=�p������1Z�g����ِ ��7^쾡�9�y��G�3f�gw6� m�h���`_3�i�2��Qx���}ᣣ"��'�P���$�◗퉩'YRK+�;g\���H��01S�H�^是�cɨ�����<	>1ļ1�yB!K�b m}!H�>�).�yԯ��XC�J����덯����vW'�6�۱s�Y� ��E(�(��~p�:�xU�VFP����������2�G�����M����?�%���VC���7������wV�d��\���ح�֙��G0.| ��,^@Q���z��SZ		�|ڡpӪT���������0D�4̠ɑ���?�W���� @�oA,�b�F=�Y��0����\r}9e+�^_��|�;�g��u��&����L6�:*/S�T�����a_��g���E��l��ѷ#�J}��G�P��Җw�{�[�i����8�l�'~ҭ�=�i��@蔈��@7ٰ�x�}1d�KҳYE�
�M��F�v��0�.�s6���7���u��o�y�r~�S�߆8�r6�(�
��ɀ��9�r���V�i��rZ�.�k��ry�ऌ�А�N�M�AҾNuc����6������I��[�sT-���1�{�UJ���i�/V.�v�zW�)�0�m���s�K)���GlzY/��"��k1�f���l��a%�\%��=Ӳe���?o�l*�9-����0Y]�z�-މ��A�-�N��Au��Ϙ��[E��Y<�7"����I!�<��/�(�V�De>�k�sF�/��%���4�H�O��5�� �(lN�������1b']vb�=��'x��Z��܊j�f)�*�)k�^��+�	7	�oxr����3X��boY�0�O��+(����RɶP��>�����H���Y}x�8����2�U����2N�Fe�:�6[�V��↔V�D��M؄��A�{�I-��	�w��x,(�4���Y��è���9���{�gT��a�e`=r��� ԛE�8g�2.��m�"}��)�NrS[Z�g��9,�f���Ĭk�R���E����Vl9]�8,������z��Q);y����an�C���*����3[^��^�`��.~B� U�ݣ����r	!�4�Ƭe��<�Zmɸ������qݰ�3�Ǟ�0��������I")��ڠMM9�lY�q����W�'��ڂ����2n�Tq���(�s�䔄�f���&}�mja!��SB�9<�X�)���rZ[�X!�P�����E-6ziP��$�]�jL�a�?~�o��|����Kmh&H�SרbN7K�^����Y�r�  ���f���!>CtЫ�l5�W���;�B+E�L<�
�(��%�eA���p���&:<��K	if�7���h�.Ag�T���h���i��?a�G{��e7��|kl���tr� A3�?���[���S��蕕2 u��Y��	#A#)2⪊�NJ4mz���D�׳�W�$�L�5i�i�VZ(d~j���N�!�
�SN�M���[_X�߸�9���w � mX��\b�H�9��Ӑ�f%.����ҵ[� ���u�B�RȽ}��g���&���7�Jh�7"����"E;�h��Y�$�s�o�M�a���J�^`ˢأ@�A��ʜ�c�`,<���rQ+�V5�e��3��ꙶ���Qś$�W);+��?�����A�S��Y��oYBq�a?r8�ܨ��J�r��u�a�ܕ,�O��1ߣX�,�sJJ���]_��5z�|������Aa`���n�K�f=���8e_5%��*�!N��b
NQp�U�n���<�0��/o������ֈ�����J@G�r��ܺ�/j/��y�����T�'z��F�>�k�Hsug {���̽��ϸ{�=�ھ� SZ;�*�����Lڐ@*M��y���ɉ���)V��A����z]��"��pY28j��m$�2UL�a���f&x�|y]Yҙ1��[һ��F�Kv�9C@��7V�TO�X�{.���;�ҟ��D���D:�M��A��c���u�7����E-�^�-���4�+���pj�S_�H�VTHi`�.W�,��!���=wO���m�X8��\U>t7|`�N#��e���5�����%��b�^�!=A��E34V�xV�R�sׁ>���;�;}WD̆.ݧ���TעJ�<��脏�t�}J3:eo�p�]��p���>�*;���d�i1��)�-��:t�k��h?�C���4M�8����&���)�$��31�_�6�n|d�Lt�Kƌ�xp�gƏ�r�ؕ��[�e�0�C�s�?�4� �q�1��i<�ߞ-��f��!9e��2u���%X�1e&����?�(@���_�z����b1ܡ��q�08-�@O��o� �^��w�=R�kihu�.����&y�Y��e��u�^9�{�Eq�.�Agq����x'? ����y�!�;��x��R�D�T��5�͗T4�f�%F��A�F]��ڼ����}��>U��<&\7-*����cҤl���Sˬ�12�vJX�5S�Q(nH��:�af*�z�	��gks2-��҂fד�Jd*�TI�I��Iۗ��8��d65���tu��!�ۭ��~�Hvx�f{�|��mf	'#Q����K��.�b��dԴ���۰F�R�px��e��u�W�%��辦2�� ,i��M�i��`������>�pbq�z���ȶ��'�s�1i���F�-D�L�V�f��I	LC��ػ /���X�%��K|��߶���K!t�7Z��]�)=�y>�JJmٔ�6@��n��(zQ��q�� z�������N9�tAv�Z�Ԝ�y��b�m6X�5V�-*�����cLW�#͆����p�|��X��g��M��^�Y</��>{xʤ*lv��f楥o�
V�Z��q��i�xJ�]D�hÚ����_�z�GEB�FG+kGd	:u�q����N��V�c^t傜�v�vU���P��Ǚg�K����`�=.�E {P�B�
`yH�V�t��=[#a�]�y��k�db�����@�iɴs���ڂ�[č*i���f�GEQ�1t	8ø\J�l�������Uǔ��hȿ3�>)[k3oR��bJ��^��D�����k��6�Cc%�C"��M�g��r��g� �=�z"��*�⤗��KS�7����\�G�'�ra������p����AV蔜���%u���ڸp���)m�kIK�R (�U#�SZv:���t)�ك�k<E�dų"�U7듦��<.mm4���U]��J؅�v�BNc����S�$��*�7�"�^�]��<M<�Q�s�Ӎ�"�JkzԓZ33��08��Sy" ���o��Cb�Ib�%�_�@��u���KS�G���dقř'�Z�2-P�}g�j��L�<v�[*��b�iiT����5cP0����c1�-ݜ�8�ĩB��&�]�������r��Ĵ�R˰��O.01�4��|N�t����"/,b9�����o3�x��  L���	[�Mސi�JQ'u�&%5qb�Aj�Єs/z��4Xu���)��X�B/��0A��� ����1f�=��ҿ���a���7���;'&d1̏#u2V���6ޭ^-�ͯ;&���(�-fBt�� �2^���:��M�����#<���x�j����a���0�1 �����u���BWh���8
B�s&	����p%�a���<�!둄�X�d&��d�ޅ��� *��G;�W	W�v���R/��9Y��S���l��`��y4:�W�~�}�^��0eK�^lO��mJ��~�,�E������#㋦9Z�>K��R�E�z?��L:$�Yw��&�qP��PtJ6]7 �3즹�B	���y,�d�A>�tX�0(P�)]�3��ӹ��{D��7ph�,��%P욙_ް����|:?���D�C�Zz����C��L�^�ʶ�,h%���(;9����Eꜷ~E� �M��P��6�P|=�;D��]h+xXL��;q]`8����F�x�ëc[a;|w��������i�����g�0�W7�_��&�qf��H�+E9����sp6�g��!lq�9�O���u��UD�Q_Ӆ�V#�B9�E\��E���
��--��s���\��߃��x��U�)�&�1�ժ��LZ6�\wu�,\9%f�6�<�gZ�z�.rI��C����/�+gy�r���eWq�y}�s�mT��aƓ������=��ɶS�/�*�8{	���&]�ly�D[;�eJ����[>0�� �<?V�aa�ۯ=�hh�>�ؖͩF1L�?���l�Q@-�Ŵ�Y��j%��^�5�Z���Y}�:b��e�V-�ȍ�+'Y�E�XZ
/��b=��Y�S��\y�����m�W�z}8�)
l��8���9l��Z%����sj[�5Ç����F����}L	����&ہq�S΋�&�G�p8�����^ B�ώ?�-�6�*0h)h���}.��[�v-$�y`�r������B+6�I[��U��Y������m�?cC�yPP#�E7ś]梑D���F�"'��2w�-��$����sq��LIҎ��g�`X�,�ৢ��D?��ʶ~�������"+S�ɛ�j͞�ʑ�6�6���v¢���������Z�����8�,᥍Z~�A�x[�����L^���n�
�1��`���n�,�v������֤�`l5��������yjt~�糗�Պv�6�2�M9�>n�+��O�MKو�)��d�g@����<�
y�5O/k�����a���Dki~*%���7Tx�#v3�ʎ�!�	��G"�4�4O�h�ǧ�kA9��ZS�G�Z4�D��#FՏ������!�1�H�d�o�3�Ծ�t��4����m�Q�>�-��̂[p:����P��u��+E�26������j���4U��ᙷ"4���,��"��6j�5g�|�t��Wпo!�f���h�?�����
.̍}g�A����Dz���MkN��������٨��@o�F������w�
�d�1�g0��G�^�zL��%Ӊr�m^��	8>^�F����cD$����o��N��7�<�dH����Z ��%���q���?�Z�z������4��� ��3�m�A�QggS�~�H9��l�؊�D�
g����6H�0�B��3����wC��G˥$@�ş?Ŀ���L���ng�'�M	��w�����B�	6~�,�����u��y`�3@#d�����+%�l� #��a��u�̐�H���G�H�^�-��c���ev���QV����-��X�f��7��U5���.��"͔����k�YaRp�Y�l�A��-���>��w�~��y[�dh������%0;��-� t��2��A6�zS+���L�̈]{D�P�xD<����56��[ɤ�	��t�HA�Nl���[�/=�8p����~�}�7���A�Mz�}�l�@5/�!%���W`���o�C�;���l5b������ֽ�Cڢ�&�~$#H�,����s���/�3˚�^w�(f޻Q?����i�/ f��0@m��]���!�1g��%A��ֽ���=�)�$4vX�G�9 *�XCqD�Ħ3d�Q�y+W�(�0�u
]R�T�땠�@jK�K*���ۺ����R��v&byJP�m�,�'�'�~	�?�6���0�A�{ϝ^ =ܫi�T�M��pZ�6��~~D�<S��&1�z�E���f"��/<Y�IYtk�Jx�;D�Q��� Ʒ�+-Ү�0mb�)B��cl����k������SN*Y��w!���)���S;[~<7������D8�#���y6Z7��P�[_F}���q0*��+
H�w�sj��D����	�)o�]$�tP�d� �mWfHNJp���ƵC[u�V�xhJp�~`���X�38�~Q.���'.ئXL*p���Yɰj�Ҳ�P�Q?�8gg�njfg��yb~�w�i{~��{�֗��`���]xs\0��Ġw%^���tؐH5�D�!ES~��+��11�ۿ����[�����V
�B-��"%<B{�V�l҂��u\�yj.��Z��B���&�-y}:5s�7I�K"�!%2��b�Q�Vsk��׆iũ���-��{�uޑ�%�/�+�������F�p��G�X�dz���%W�L�C�d�u���-ݼ�.�*@�\�ѡK��ׂ\�cJ��Ū���;�8d�J�Y����8�M���1��)�0N�&��	{���7vL+��N�6XDxK������i����S���З׊��U�9r3�ϩ�h4�i$f���M�� g̤;B��bc@�)��Fnꇲ=��M ���l$!�}>+�{�^�~:y�%� �sR!#<�B��b��|L��c��œ`m,I��*}^�x��M��hT��0ӽ��fb�Z��58}�D�4�F�7^�Qg��RB-��V8�"��� #�xe}���	��Kެ>�=~ٮ��'�`�q�8}���vNݰ�u5od�˕�wϐ�+�}	����v��׼Hn�\vyL�zAC���H�&��<07�`S=am��[z@����W��j]�x�R?
g;]��U��~���
(����de1���X���)::�����AF^)�4II�OC���ٗ*Q�5Q���?�=��u����;�Ē���qڢg�}Hr_��j��U�6�v�Y�*�Q���ly�"���I5G�E��J!�n�~�1�t���rǇ�>M1[*�78������4ϩo��m)t�K�ct�̈́X���|�c
�1.%�����YnH�u�Tq�veƏ��R������[�6��:��UwN��d���x���VЙ-�6�ڇ�ױr�0�e��񦸿�Dh�ti������nh*$�l����@� 8*�^ԾV�(�gk���r3
��np�DhI���jU�e�?O6���-� N洝b�T���~��*"�m�>���\���ћP�1���Q����"{��t0p�P�R�'�d��ٲχ�
,�����:�����$��ԇG.d>m��0S1��|̞S��H�J�j����R�o��XK'paV\뾿�n,�*hx�sw?�����*�g���<�
8G0��e=z"��a�_mf�2�$��5No돞AC,Zvt8?���k��Ip��M����WM��{�� _�u!H��&R~��'�#�VA�ijM,�����ۗ���jBG�V]��&��g���Ƚi]t�R�)Jv����!����`"�q�O-^^;pp��@����*�N�.�/P���'E�?��E�]J�|��@��v�|x��m�P�Z�r����D7�A����h�Op�Ac��1�i�I>T{7`�'�����3�A�7���'
|Oc΍�|��CU�7���X����p��;�Q��!q	�F�[+�|uJ/�hܚo4Z���?�O��a�߿�.���j�Z�����֟�����@6�e!A���;�7�6�g�=�7A@��n9Z����㨽z�pVd��O�X7g{�	���tt�+�u�\�̝���jK�1ٞ��MVSV/��"��=����i+],��6�1�[��i�4��> "�MlEI��V�@��+�T�4�1����M�������Hm�,��o�����&૭��D�_%|-�;����2[l0ww0��X�������.�G�����\A(�AS�f�΃��G�Fq6f7rx�΄y�L�Y��4Q�؋5��͹�B�vި���`k��3����;.ݰ<*]3&�ۏ�wʩ*sirAa���P�D�W�4��&�V�F���,S�I\�1-:��+\�Lp�������,$�����C����g�}�9�O��6!��:,�X�u`�<sߔdw��1A�H���x�������kA���51+�7�Š�W"9z��z�M��G��)�~+�-w
�{��o�z�e�|ō�l|����bz|2�A期�Lid� �xK3MP�S�r�������(mC>&z=<j�"c��=X�Ӳa� ��}�ف�#�V{Y�_;o�uQ�6���b�Od��Zq�C-�����w��VmM��-���,���DP���l0���(j�0v��15)�^�X(��P���� ��{}�,U������i؍B��N-w���t�D[�K$���^�ۧ�̳�K��
ؚo.`� ���Z9�@J�IH�EJ5�_��}ͅe��M��K�'j7w�^k]Z�p%�J7�/]n�)�¶ז=�2��_Ρ�r�����џZ��S��<2����k
�����Q�X��t�S���:�"�6�y���|S�Ȭ��ҕṄ*����� ���7;�}��Ce2���w.�2�pۘ��M�u18q$��s�[g�Q���WL�>B�<}�`�R��]��l��D��Ui���fQ�n�z�^.B�[����9��n,3�BG���뒴���ݢ�Q����
RMM"��na�L�aHjT�H���j@$M9�(�,��:*0����c��� ��F�"��ng V�q���-����,'�\�4ge��QL�?��8��EN;*"'�hA�	��fP�0�Vג($���c��P_�2�\�bv����emG��#C�`+-�)�V9�*E�G���*���``*u��T�S	���}�HU��a�a6`�8�A@�Ь�5B;p\>_�-�Ħ�LJ#�:�m]}��Vَ��eH����v��1b#���f���� �bu��+w$�'�a}-�8�3�+Nn�%��pLE�G�*6��
f��X�
�����%�(��a�b��ԙ����DGxD�)B�L$���Շ[��b*����c�E��YYZ�
r"��O���WUO��Gb˔k��
d�5ŨK���p�5�^��V9�Er>�t�r�e:�O�5�Rq�'�㶯)�WP:���iRGO�Y�ڡ�UP ����%�E�DP8�q���.���z-��#2켬h�/���ZI�I�n5�zs���M|��R����5��n�AY�M���J��Q8
{⻫�[����&9����H�$�Qc���;��6��q��/�P�mP̮�d�V��G؍#ә�V	�q�HN����Jb�f^f��8�G٤ ��k^̲�4"��,?k۠��0���l�j��Ӳze���6�Y�	{tY��4�4Ȧ���LwB��b���z3O���;�1�Gn){�����'r��i�Y��I�(ː���!R��O�:��4-��L����uS�>رp�\`��a���u��K����0�ֶߠ�P��6��֤��s rӴ�C���n�G��c ����/�:�;���c��\~�9��<�sd�1#��k�v}�[;k�:5͢\ާ�_�J��4��h��xt�����Ȍ�����v�-#�aQ��L|>8AGN�쩼k����^vj��1�m�R�Qk+�U���=u �ّf�?v�u�Yٳ�HmA��b��G���զ-��􌱌�0��%�5��.<�W��?�DVw��M5�I�%ώ/rߨ̿���z^,ӎ.߮u:�H}���p��5;��T`,��Җ�;T�pt��[���4|ڞu�fн��p<�rO�U���Y��MeE~�>]�`��	��ʆ��m�4$Ը�I'yrS����p���=�G{��b@���SM6��
�d�dQ
�ү���U0���U���s�W��� Z����Q�8=3j߅��+ i, �DĠ0�i��NLO.�q��񡤦�+���W.4d�LZڿ�C��1Fv�!����q[aG~��Y��ʰQD �a(S�Pm��~f�]��`~�X��:<�(3�j�v�p���\ƹ������3s[��ŧ1����m2�S�!�O�-�>�8t��8ב^f7���09��㯝� ���b"jh���m�YugO5�\��_�@�P
�1�{l�<ZŌD�EX�g�A,ۑ���B�>Lt=���u(b�_a�h�箌��F�e��up�'2��G��:2�|1� YK��#��~�Jِ󕴬��j*��֏��i-�&�\��dH���ZՄ�5er�rj����r�ܹ
�sUZ3�7K���l̬�y���v�U7�r��Iw��H���w�I�/�����Q�U���ˆ@�o%�r���R�8&d�w���0� �KC0���=GS2�4����w^����&�����\(���ڋ�����KP^N@)!����%f ��j@,�������7��=?$h�������)r!��K*w���8�b'o��z�fN��--�!Ҁ�NF�l�vre����L��]�ubv2���)��K8�'v������xn����p^P,��N�XmŲ��yUۨ�=�*�=�H�m�N�x4�'�\��x�?@��˹���4?h�BʿF�� �$������E�c�!e[1��g��K���DĐ�;���|��%Ӑ]�z�QJv�jZ�U�c+d���跰�襝qH�Cv�\�,@(`�&�Re���v!;,���s׮j.�4i�p��D�ފ�Hsg[w�'�����ժ�_���9�$5��7�w@��mZt j�:~0\�ߟr�A�~����0K?���s�A@	1-/�<ē/*� �^^N_HgG@��R�7��&�rI/%�<�7��=O�U u[�I�����G���>x���UM����sZa�b������I�L��پ�*KIߣ�=�BS��X=��A��+�{�g�gki��Zwb'�ݰ��H�a��h��T'v�bAٟ�!=���و�
�D]:+♉�Ї_z{7bl�93ˉ���d�^�<��)z�h�V>y_�����K^���ʄ<6���� ��[6Ɇ嬬�1�@���!���m�)���5n�tRt��~֪\��dR�@n҄a.�U]l��H������CP�F��J�cǶ�[R�L�Ń)R��;"P��bay y�A�e�� ���T?h�o9�#��؏K{U�(i�s+�:'�hn� �w�����@���y�>�$�X�yZj>6�_O��>���G|*$��}����/U�v�7�.��'ݡ�u�@�s���9��Sت�{-Wd�C��,
^�]?s�gNW��4�6R������
�!���� ގ�X��%��3����3��A�T�h���~zVhŰi��Zo�	]g\
�U۲�t�ʒ�S��N�G({�n0����.��Eb�t#�A!f"�'j>�q�{ ��;�]���p<��e!�[:��F�q���5'OW�/�HЯ�^��p��-�Jam�������y�'͸��5]F�_��yt���>�	�A`۟Fi���y�&����������~�?�o#�����/)��Ke:�\F�9�ȋN�j�*�y"Av��k�Me&�z�	_�G��@|���W1ڌY�*x��$��.O�yh�k���$��	���8�v�<}rz8oM�Жq){�F� s�w�c8��z>�o�q�o\�C��0��B�J��嬊�r9�YQ�>�(�$��"�ܬ�ؐF�ݱ^4E�Y�UΊ��=)�,��o3����7�SmWc�;�?C����z��g�P��Ly�X�}�%^f�4՜��Z6��a�=��J�L<���Oē�mW�Ĩ M��ru��H�/�{C��}�g-
�B��hT�c4f2��d����=�/�f�`Eyd�P�B�(z� ��x�z���<�������zn	s?�o����Yd� �j��7�V^hW�yoE=�1���|��ӛ�-<r4��ã��k6
x���Cja�Q�����,L�c�uW���8�E�6��g���n��LQf�.�Ubp��u�RhO���c0�@���S�N������Ҡ17'�q��@�-{�^��k���a�*��p���Mm��`̍���Y˹���Ő��8@ ����aԐ��ٓ��4z��ح���Ov*�z���x��v������w~#)	��W����j���$^���Սރ�lG<���/<���OJ/32�(�!��ne�M��q1l֞�
�c���x�� Nl[Ϊ⦀B֤BZ�$eԀl׏���P�����v���^ ��b��d��S*�w}
Z�� �݃W'>�7���7������<h�VS�X������Ń�o����TK�L�����e$�ɛ�0.��Qqs=���*K�{�t�����g.hT/&KH��Z��w�@0��(��j�Jr4�_����T�#�	o���.Dj�\��n�4����]dW[]�w"FzZ7�[&�c���Y0��՛$�i���C�1��c;P�~h�����3�c�&6/\5���%E�8��M��u�L\<rXif�A���Ks�"� ��:8Ćҷ,�Xbr"N"���p5^�J��~<o4��V[Zb��y1��}2��a�H�r;��Z�ͽF�"U0d��9s��5�
���Hv��<B*u�#�y���"��� ��i	�R��pJd����P�"�4�FD�z��y�7����u���C�>�xS!Ǫ�+��x��Hv'���-#��\����M�T�z:����Z��9<�b���	��;oDؙx|ߗ�E/�V�$y�Gd���1eH��1�Sh���ёc��򎎶H�=�$mpP�V��e����F��j�K��~��B���۬,d#��eA��VJ�iC��7�[�o9�� ��7���R��[�8b\z�B�����K�q�{Q��������4K�	k�&ԛ(�WUAv(����mU�y!{�?w[h}�M�d�=�x��]=	b;�A~t%��9 �6�W������œ0�%����vxS7껇���C���f��� �,F_%�s�罜<��o�i�v���?V��͈���C�Y�u���T49zgd�C���7�аZ}�&����o.�����Q�I��7�G0���z 5SE�h1!�o�;�椻����C*q�Q	n���Y>'�(�cF?�r�=��� hg;b�~��q3�
�"+�խ1e��Z>k���:_�&#x�2�@���`V�}��XRm��ݍy�΅N8zvĵ�'���(V:�+�8��L��H�Y�	�� n܎�vr^8Epv�B%�'�kΨ����N�v�_�ҡorV.��T%|��R%C�9�%P}���S�����
/��-�K��B�J��9��,G"��r֨h�r8||oo_��	i����u���(��~�X�zԓ�>�\@9	���(�ʋҒ�e�������	"3�W
ߋ�s`�~�<��z��$1���v8*��ZO�f�\6�F^����(���GFO�,�PD�;
�@��z���Ɇ�I"�������lB�JQ��E�tі���K-�ʾ�xP���w׫�����/.[>?MXP�Jۂ�.[_�r�P�������VϪQ�<<���1�Y!Y�}��s�!0܈��͏�1-�/H���M�m��1��Od��ݵ	Y�+�>Ϧ1�����W��֘�G�_��0n�9a꘽��[{�u���9I���L��-u���_ϸ\�	*@�i�^b��N���X(S���A�U#��,�/K���V�r���RAЖM�$���T�:*��]T�/T�r~a�H(%�WNv���&ָ���o2�N�]����W����,}���y����LH�G��iz����c�܊�9+���r�����0g+FX\K��8VT��o!�!�j���`>	� F�Sl����܆F���I��EYM�i �>w�,R���� �%�B���'B�['�o���΀��ZU ��Nb4�&��+�t|�f�&�������GHх�Ln����7���!sl��f=*���H�0O�0y���A?��\8P1�Nsi;
��w����s�������������B���#M� Y��^Ay]�3dY�jL��#�01$d��_�z�m�<W:�I\b̳/�>O8�⊀����jM���s��c�-��#�15��1cҚW������8��Ƞ_A��&�k
c�(k�!�{W�/��,Oı�K}O�d�*��R�`�J��#���/mT`�8 �����1;]��L=�����Re��޸"��m�\	J+���۶Jy����:�,wD��DР����� �������.�|�'����R�Zs�7���1z��{�c5���8��p� R�&�bӥ�O���͔ر���2�I#�PlHt@�H�d�&�A���M�����:�@SG�XH���#�{�Ǥ�����V�,}čvlN-�x�V/J<��l�?��6<�iKQ�����H?��G��ϸm�D��UO(�&�gK�"�=��;q�u5"�u6wu�e�K��VzWpC�ο�!���Јr�[�=p�3�y&5l���X���Q��j�n�Ad�Y�8�F2��J�U��
�b�?����k�j�H����Hx�^e��ޔi�� ��ˀ`�{���A��+�]�M@Wg|�s~�Qw-�����}L�6Y���٠��w�P���S��]����W�V����0:}�	:u҉i�ҷS�&NրёƋU����"��bU��]޻���1�^&���/P���p�w�33�?�s�"���IB�q���z��:EX^5	�n1��µhq�+�[j��D���0�,T'�\
ݰ��OtɪnLH~�/�2z�:����k��hA�V�q�ڭbP�^���e@HB�9�km���LGtU� �1��x��A2.t�7)j����n�cS�&˞cNc�3�B���^9B�M���j��c."ENa^FЖU��$���Z��Y	&�<c����Q�pu\�b������l�&E�K��PV�&s]��)S���[)G��������_(�����f0��Ư�-���ۡx�<�1�|��D7����Ig@73�ק�}f����#�ގ2��5
!٫:\l��}P+)���I�<�`�=�	��@�4 ��4��յ!i�q'z:��8�ofخ��!�H�P�2�4��J����d_��Z�f���6�v���e�^�J��&oN�k�s�N��y���//v7��g{t��� ��*I� ��+�<���ec��̄��� vҬ��^ ����Y�.�k�ZGS2_�윦���rA��اP��j�?4�	�`��O��B;g,�Q�b�2�ƀY���m8�'�nl��;�dx�';Iv@��C���!Ee#R�����i�w[xg\�9E\1�J+�l��XM����	�	g,5qW[jőD��g�������o�4��~��S��m �~P�!�2~�ֵ�ު⤕lO��&��L�B{���}���#���C���m�v<Sg�����]͂��V�����BD�怘�NV`���f/�B�3�`�*|W^��S�_��	G���/7-ěaNCA&�2՟���ץ[K���h5�1���ad��&݅8mq��Mk_Sn��۹��.В����� S��-��Ĺ�
m����<w�td�+d���*�]VN�/�Ktr���N>[@U�v�f��6�};�qC*�c�)��_Q���&�y�-}!��B�>^B���\-����ʬ���p���E�f��=ua��)�|X�HC͜� ��U�������H�*E����|��V����s�R������ë6�gcS��P�Q�Z�A�s���h�0N*Ȩ�;u��J[�J�k�P��-!%�^N?���������Jw��^�`j��=O������l�p�ڞ�߲�v
�}+![�l?�YV���McfJ�N8�� Me��8�0�$s��=� ����v_�m��>SJ""Gc�K��S�����y�m�{�n��6����M;"�J�{���Je=W����0us���ݞ���������l�u吟!��B�5P����DhrҲ%	u��^�X���h��f���R�̹�����Bx��L��}#֭CVI
��{�|1�l�ӯdM+�00�g2�qm���m�j�hq3V?�
{ �� �[}���k5"�V委�0}O-K�2��[-�_ �w��`�Z����jX��0D���:��B�L�Gd�W���/��E�n���*v���%���ͅ�#7jp��V��ħ�>$�4zJg-��vi���Q`e?����~�
�
�Rm�h �u�_��Clc�6O�����I��#��3.���ݛ9��@�������딇+�G�=�=�*�]��f��>��FO���w9�	�!'z���97=!�g�Oׅ[羝#Ѐ����X��iPZ�C˺O���ܣ�xL�۔e��� .6�Nw��u�7�o9,)x�i�|%����Ʃ��7�ʡ�Ab|��أ����������F���"�}7O�?��2��M�7��)��w���HQ�H��ws�.3�S�E�}O��ZB̆������8��0��poii,�'W�!ɛl�eu�T���Jn��ߌ�1��c�+L���=*Q���[9��C��[�c� �#6��E��u��]�}d,���������J(�����X���\�,���dKXz@��Av~����],�(_0�Et����F�	�0!Z6a �+�O�C���0��#GoFd��r��y����QZ{�9"�{?�Z���D��1�1D���O�R�f<�?n3�4!r�a	����3���c��Om#e�9z���������v=����=�p[H�l���^��8�|9�/���U���6��4��N�.~���F*�e��`e%���bp���P5��MQOOg0�������w�a�&�eOvG8��U��{Y�g���]�V�L��������ԗ6Y��B�mR��-�����i�k�|	p)
D��6����\�sK���E�u�Q/�w'|!�|�S��|	=CSKaD��uV���4X��5�5���X�h�e4;\�����YW~�#�
�>����VK3�G/E�~A���5*<r��iS���K�>����R��k�*{��0���~ӇIrs�A0��P��3���R�(�:تϞ�8�]w�y���@�T3�Fh�7%dK��C;�Q��f!�,`��(�P-��{w��5?��ʋ�2��t�,e7L�|+�)���Y7/ ����\�p���:�ȹ(���#�,����Ax�>!�>�h3�`}��s
U���,���\�����TD)�D~7��C�Tm(�SM �D���;d�Ԍ�j&Xj�/f�"�������*ep�V�x�M΄pB�X�ܜOX�@��k��~�6y���].���7�{ΊϺw.���[ގ>�� !�DZi*B9�z��J��A�C�-� {DV*� )���ω���L�Rѷt��X���鳯
N���$8�
N�iCzxD	�n�v���e7$RP�|p+9��$}�&���f�dV��y���o\�#�; `��=�8pZԡ��4c�_V����!C��i�%9դ{
�(��T���Ns�Z��o3H �E�v���c4�_�<0�=�])(�LlXA��Ic4!n!-
�0��T��^�FC\?�R��L)-ص�*�/�[�i�|+D[��Q�JK�^��������`5���w�ѵ#ً�`�1ZU�#�ǈ{�*.�L��r��Y;��L˳�U7&GN�1����`'�~��|�[�y����7�ٗ>ޚ�K��^�B��B�/�5/B���l0�e�޴��g�bz�練�@:m]H���� �[Ji ;����Nշ�hv�\Р�=	u�׼68B6�Z�.R�DLEe�L?1��aa4ַ����q�o����bE�����x!�i�?�ߣF��@�Nb+��"z?פ̛��h���8�O0z����y�1���${��r�0�����[N�+��g�O��#�c"G���5��5��g�F"R#���l��xT`��4/o�=�Bp����7Ѐ��v"b�{U�H����C�N�����@xbhyS뿧Ӵ�K^Y�{D��V8��
V��)jާ�7��=�V)����L������������м��F����ԁ� �����ٜ�L��?�'u% H�WH�N^A��O���f������y
��k>Oo�����۪��{��ׂ�&��l8��61���TF:�����%�{�t����=� B���?޺����4�7n���Ǿ�p_PkMr�����G9z�Y�<�C�Z&Рت4�u���"Ԁ�3�J:K�M�N���k�/=A��\��G2��3
�b_]ѫ���+�|��p,X�����?�:���rh��z�o�E�yAv���x޽kǑT�{��N����^(���%#���)�	o}q]˷Zs���)R���A�7�r�S�#e��� ��)m��r�+�]F�������,����]��G�#����ۘo�Q�Y"ܛS�&�;�y���'�qU�5��^�)3i�?����7�,��q̎p��[��He"��z`�T*5�}=��B҈���Ug@j���ڤ����%�qR?��U�#�����S��L��x��u�Z�A�=�F�&�U'�+�k���7�y���U(
f����g�����52z�����iC�|���z��3��9�62�Wn�eo�F����p�	g�А�.c�y+��E2�N��H�m8[b+�5o
ժuiyZ������X<�2�S�r-V��[%�#���N��1sd.ԛH@8�ݡ�i�_s0B m֋B=-!��kd���+�&�����b6�����8�}`��d�;�(%�O0��9� ������B<2T&%ii>~Vߍ�+���f��Еo����}�i.77#���X�H�(/D�o�����vl?�pYDKjM�>�>{a{c���E��c�6Ź��C��3�;*������RH#_T�̘�W0���YL{�8��X�N'Zh<�3"A�j{���hn������
�I�����_�s-���X��G[���� Ps4��0��0{��t)���O²��tȘ��3��Z��"d5Y��ۉX���o��!QqN���H}w�=Bc�Y[�yw9�Ab��������e�48�Ҡ'��0U?�8̔O�3���&�,L�����8u�{ļ���Ǫ�=��,\`�lݰ��S����O�l�|�I��W�l��`�n�W�{0^�.�$dq���ǘ�d�E U ���"r��W�g�[+�A�=��`0p�(<������Ǧ�#��SE����$*�z��yio��ycM�נ��B��W�)j�Q&����3C߀&����$�Ѥ�\n��}���,Ȅ���)P�M�%$�#8���I�aZ�Vý�DanL8M��Ϭ��f녉����u�4��J�A2��"j���jF9l�y��bJ��Kt��@s�V��Jӓ���{u=(#�Ҁc/��E_���t6i޽Y�!�7Ya���=_pW:'����x{�4O8�ʠI~N��p_�d�B���eMlfyH�@_�`_X#�G���UTX�5�4�ˑ'�w��aa[���4#�0g��߷��M�H�pr��fʮe�-S�x��Ә��H�ad�7�.R�

�߅�?>LCh[�jۖ�$���r�����!f�l�d���*~r��|�k��,���N
�����./�Է�K3o�T
�H�g"obKeɠ 2��~����v������e&�|)}2]"���E�2�G�������=,��ֆ�� l��4i�d�s��4�nM�Z�H��3�Ђ��Xh���Y�R8wx6������}�P�f>��c�*{O�e��; �f.�9���,r��&�w�>;�R^��\*,���G7����)�*cJ`oP�}8�N�ܯ�$�ZE��pv2�������`��I��`U$���05|��I�b/�驮V�.*�+�IR�ݜ� {��UMu�9���M�^<ϕ�h��BZ*�<��c�j�y~�OE�'��N��<�i�yϘ�WGv7���gH:�O�ˏ�'��K�������3�v҉�R���ǐ��ڸ�-4F�J����i:S@���Z�r��,݋Ǹ7�m慍o�3#$�%͜nӣ/ٿ��1z�����Sk1VW�{R�K��q�{:Y�S�~s�\���+6X�E�����z�}���)l�2�(��Im���5q���E�Tr	aمNAt��4!&%�{Pܺ��n���~�
&Gx�T�7�\ki��xy��J��ew��� ���Ry�H���Z7��~c��;���OnO`�l�T�T;Z��t�=�%D�r+���Ot���:�j}�c)�YO�Hy�B�=1uN�.�0/o�4�>kJN{]�Q\��v78��_!�F%g�E7 i(��H*#%̗Զ<(񷟕�i��x����~"]�։��,��W���e.ƅ��֢�Er��{���b�#^�=oW/��c;^��Y8���I��-�Z��*Cf�zJ�ë8;zgtu� ��%�WESɯ���,̫�c)�L�ͅDCӞ?x3�ݯaO�L�v�Ƣ�j�Uh�ڇ�n�i)�Љ�3���v��r�����kG�oi��I|�[Z<BD�#��@���:S���$>�5�N�7�S���]tz!c娄�Q�N��yC�|�㸋?��x�AX�1����(
k�, 3���0�E�� �;x��^u{��?֎j�oE (�A���9�4�H��!�� ;6�� �xu�ثי���{�Ez3�j���:o�J���ۖI���ݦ��0�qT(���F#R�	&.5�#�3�� ��F��!�-�fk�ga�G����53��fJ��o;��lr���� G7D�,lb��A���@��O@��������8�n4��:��u�
�rV�~z�X�,��A�W�;9{�|��I%ɗ}��߸�0�ǜ{�B)/-��*��C�����j�n���
����p*?���V6:��G�&�]d�O�z�߷��[H,OAzS{�픮1 ���S-֡eR�E�ذ���o�A�h^"@�O �ʓ�<��,[M�(���%�p��3}^�݂�Q��	(�΀�4h��� ��ŵ�t���z~)9@��x��|��[N`Z!R"P�Ă�n�-��о�~U���r�A'8̔�!{E
8��\2=*^��Ĳ�:r54�t�����~���W��zs�r�����h��6�Bl�N9cpc6�f�٨��r�G�1=�1��hڜ�}�U7�!�p��K(-��԰��8$F@���m�[+5j��w0(>������9e�ؕ[��L�ݥ[�����t�5;4H-~�:b����j�b���H����2rR��������nd@e��V�c���_ZfLJ��E�:�I>����3������~�*&���H�\8����ne�+4�~ݟ���u��+��,\�P�Rb-���rQ�oz����ף��"� ��C�2Vj䶔���D���^�bL�B�T>�3���{��u�h����������ض�<�Ҝg���
�,徻��v�ᑜ([�a�RDpO��ƈ����Hp��j9�fJ<ꖹ�s�����M��������5�Cڥ�	Nw����(����\:��o�GK�hB%M/�F� B�-���u"�V�g!\��Z�%{2���/ ;	�U��b���K�{Du�Ɗ�Y3�`\Nf"�<Ȇ��Ko��]-�Xp�b�>H�*"9P#́m���Cסb���K�u���4W�����l�	Dc��6��\$C �!��T��@����}����5�����)�`����x�Ů]9�ǲ� ��m�~��\R$�_���
q���ѓ/|%}/y/�؈�����z�%)��D�>E�ֆI����v7wjs�b^S·M��nԔ)�-@'�I��1��U�*�� �F�/}�/�I�h��E�(�㩒��iu�w�}�7>W}�X�<.��~��1�8~�y��9 �+��$5���l�ML��-��<���[��J����ܔ���P6�1�:���=�c�/�5��=i�3�����^�X�t�0IJ�Ts�`hΩ.�$a\$�͡����q��%�Ȏ	ݲ�{�\GR1ɱ7&���`�mߋ�n8� �MF\�F�Ͽ��� 6�[���\M���;~��Ǖl�=:�&��+�ݢ�nf��3��+gBCo(hX�)��q�'��;Q���i_5���5��OSnĚ��*�F�r�@�&ڧ�b~0�[���&3��L���k�� ��N��}�OP"�c�ﻔ�_�D����v8Ki[�fGf��<��I|4�>P�i���+DD%X�t���d�}��ߝ�⒀G�m��f#l�.\�P+�NJd\3mZ��E*e�>Au�.�����F�%;u��췂�N�ϻ�cޤ�̳�8C�+��'+�؃��w�&�>^�ߜMd�FO,a��l�j(I���!B �v��A�����_D^=Q�y�.��\Ƈ����hDb�0�G�	eɓj����!G.�D�d��d]��Ӗ�?�������k5l"���= %��V[�[ˇ`��A�$p��	���KFed�K�X�N�����Ѿ���o4�s{��]S!fٓ���&�,�[�9�����約d����*��ø�j�,93ܚ|7�����7.�S5ąe�Z(��E٧�k��
��R�S)�=�up����"�${)�`� x��k����ﱥ?����˚ݱ��F�hР�c�F� ���7������mK�ܯ����c�����3�м!qa��Ȃ�t���=�@�6v����)�26����d��`�%,<��NX�pGz�A�F��v�ԧ��q��wt�����+��BD2�e;�G�=}]��O�=]U�޺��wZ�z����r�u��"oc��{!1b��a�,��6rQp�l�uq|q-3�o�NS�H�EI�?B(���@!��d�]q�U@L^�_|�A�V��XR�0k9f�ÊW�k<�j-$�o�.@�L����x�z���A1����x��qN�9R�LY+��w1��!�l��m�vUH` �F;���� >%�|�m�|��_�U��R�������Cs�&?)��������
��rD�����߅j�d��r�2���XV�������gA �Nw�K��E_ӈ�u�z�{�<������lw�Q_Is���1r�)�S:��CZ{9�L����$s�L�s�Ż3FfFL��.i�,CA��|�7����C���.c^{�ᤈ�IIp�P_��|�Yo�{��"�����!���w�����(HE�IP�o 'LӲ�v�l�A>�bЧ���Vi�G������h��.����f�11�� ę�#���FD��U!�`�Eح�T��~�v\�<-�� ��9)��v���W�s �P��5/[�FX>:�hp��`j��gL�MA���$-�R�CX�R�0�w�py�h�ɷBU�[��C䬡y8&�o_��O�}��\���>nt17lv0	oe?{eql%"�"��d�_�zw}L%���M�lZF0ެ��*9�`��h��Bj��N�*P��^�w'��b��`�L�<�Vj�k�DE��s$�CW��-���⢂٣�z��M���^B�b�U�����?~�XU�G�o��1�=���0� �`{�=��O\��^��
��ON��`�� �sA@QG{u��ɻh���E�?�o���nڥ@#��O�.=�r*`̵��y���1Y6"�f�C�[��a��eB�+�:ks�t}��T�Ҧ+Lk�W�MP��j[�̦�ՉCDBi��)v�[�پ�6�5�w����7 ňUo�EU y�Kz�4�`��ɷxP?<�ʟsr�����$�뉀�1x�;Nht>�������Ee�{ב�S��
h@Ǒ)���M��]�wrP��a���''��a�� o��j�_��!����G�ˢ����x�$R�Q�����z��O��/�yR��l>y��_��N��렟E�K�LjBM�*�z���t �Q�d���O�eMG�B���toL�ڕ�:w@v{��	�@8p�=,�z�ʦ7�}H־�@��A�Dx^�� #uC{�KU�bc@����c�oO�ܥ���ˀp�OPa�i�d �B�ftpU��.yO���1�o�ܧfr�ìL���
���NJ��)).-t���7L���B�7�\��+��<,��3 �]%-��Ixg�W��B㩷�n[I���L�i�8�M�0��窄!'_���,Ku�>�#PQ�;��r�02$Z�xV�h���˓�i��i�
~!�J���0Hr�E�.4�w��I��_����<�b4$��h4��t��{�C���{�
��j4���uj����9���������e���7
"e�'<0v�8��A�������{�mּ��'�+��/�r륅\���.4H4ǀ1@��86k�kaF��lxY|
���ǳ������_7������h�J^r�����)3���'��۝	1E쑆P��Yr�곉U�n<���t�bj�Z9F�E%p����[����l:�@+��� �B����CT���8��Ż�v����{��֭��85�N�����E�������FG�y[#�H'�������������a0`bNE�(,.��:��R�צ�!x�b�F7�j�K|}��-��x��ӯ�.P�@�}�%!Y��4�CQ��d��+b~o]�{l���
��[��#e+	3���룆\�\Za�`�4_C�ѯ��������-����djP�(,5���US�b>�x<�jV8�s�O��܃��gԍ��Δ)��i�l�˹�d��(�ͅЎ§��]�la 8~��̷R[������Z�En{�o�k0P|S�- ��F��]z"$��e�k�'l����O����hu�ǤJxŠ�zj�tt�^�u��I���|��㹺S��R�֌��{@Ȑ`J3�����'�`�ޮ���+8�}�{^*���ͤS�O4��h*��P��CrL�)��&��܈�&3FO5.��`�ԑ�Ԗ�@"�	�����w|4�'�86̪�i�G����R���Æ8�q#�~Z��Q"������W�;k䘍3f	�-G	��������'JV9x�He���h�-��f:�WK6��Zy��d�d��9�ͅ�'0Z4XV�L��6���n��������eڀ=pk͹jF@��(FXJ0��E��f���%t'n���(*��1�w��i�c��[��3��������i�\��m�����������,|ŭj��6\�Qx#!.p��S]L�ʖ C�#����$D�b�:%<��=	g�n�1u�F���1J�u_A���#�F��I_�#6�����Y�=�S�_~�R.��_"҆	�x���T�Sd���LdCNx�����cM]��d~I��[�c�*4��ha��z�m���&i��MOH����2���s'�tfU@�T�F���A���R���{U�,:� �y��@���p��F���,%�Oe%l��Qʥ��;?�t|8�X#Tp{��Y�uK��j֖X�[��1��F�3&�˨�oԏ��E"	4:�בo�:I��CD������S&�dY/��&]ˈ�����&`�Z����<Mq���t��JU��ݚ·�$�*���%,aB����7o�;o�.4��Ч�[��U�-���9�<��C�?��j����QJW�B�4Χ�|����'���V��w��)iW��GO��wO!��*j{d���3��ڢ�����+�+ǔ�R**�ĵ�ʏ�+$���)��� ¢1����1�K/᷼3/�~���eSp�kŘ��!��=~xz�&B�x��u��R�]�N[�]��Kd[���[E�����a$�-�����gG6YB��0A�Q:Z%?�QOM����n���WZ� wX_PS���4Uk�P����ϴ3�[\��� �1�T2���)�Ėl��]����Y�����*<`�+)���� `'m/��FM8���֟��k�A�	䊄�7X?�@I�R7�_�w������<��hۚ�aj��Dڈ�'iP�'�`@ ��]q2���V�FēZ��ݩz[����Zr+S��n�VQ$E�Шz_�n�0�n^�B�hZ��	hQ��[^��Ez�|��i�A������_c�c����5�cD���6���rf����MrǻI�{/"�>X�9�VV$!E�F2����sp��@D���1|�7">R�T��[�k�6�=D�>D��0�A���h�yo{q����	�/���o���?J=ǩ=)W��rm��"�Q��M/}�-)���|��zK�9�q��M�oV�Ԛ<nW,!��..b�[us�deU���X��w�S�����m�Q��1��&6aQ�B�a~g�tO��SP ^�����'���9R!??-~_E���m#k
�|q�� hG.�j<-hzTk-�`�+��gcj�<W#�ǻ:l7�~./�r�����dw?~"��K(��4�e���/ |8�)��V0K���􎡿7Z���g�S{�u�U�T{�$���JP{+Q$|@���<=Z=�����\'�~�!��n�����������b���
2F��&"O+�������y?Ҁ��0�"�����@��3��\m<��E�57P�켟���)�$� 2+'�,|G>��v��-T��#	�4�-|JYFD���g1�=d��6In��r���nf��邭&�,��SW�9�T�m/P�I������D�ؙx�|F���u�e`�v/��0!>��!;��0����`	Cw��[�H��J;\�@5���x.�^�6:E�s���$4�ʛ-���ڗ�R[f�l���R=ޑH�)�(u�N	>�'�		�!|1��4�g٭	�Ex�ʲ��\��<1Z�Ә�8��=E�S�i�b r��0���������o�	ֺN��ح�4XJ9����Hf~L���ހ{�g�y��J���w8ǉ��(�W{�l^���MċX�N~��U�4d"Һa�v��w�B�WxR��(���:nLְ���=�b�o㡊ؑ?�rl�B���qԉ�&S�R�+��s��9�����ǁE6�PɄG({��ܫ��]��S��+��>z�%2�hNm5ҚDS}�<�4��[��`��!*�*2���O�	�-:���pV&"?�2a�w��|Ӧ-$؁=΀m�IHά�oA:��2���#C����@�E��yhFPu<8��[�M�>I�*}Qnh7.L"|�C��7�ge����o�wӸU��Q<j5t�@?���5��73[&� �3;�V�)T4n	ބ�2��ɍ����.�a��(�����}�}]xG4c�P�>:#��=DS��V0�^�=�s0��4{��i}U�U��A�T�T�7��������3T�:�18��c�^��~{�I�2[�O�aB���K
���=��EZM�� E�� ��XQ�|��F��K�:~�(�cf@�xbN�����Caf&�pv`��h(��G��+mO=X���/��Z2	I��pC�*�<f/ͥ�v�N��Jn��;�F�{\�������]�X6ۧ
[b����/���ؐ�	0bɜg�[x�r1�D�(�� ���vQp�_�I�%p��UMk��c�*���ߘ�v.]�8{Ԡ�T���E�����E�<�_�^��Y�HOCj ^���N�^��KM2�, ��4L4�3�ѐ�jH�Ke�tH%"悔�TNp��-���9�t[�i�b6�����Z����ґtdu���`�b�,�S�r�ZW�_u�dy�����?r%^g�+�Xwb.�JMq�"26 ��F��|I�Q	�U��Lx��=L ߥ�C�h�=��sq���y����z�Mo"&?���|++Ec����f_4i� �gux����?jCǨ�6�F��W���KSE���12^��wjx�F-LDu�Q�k!�z�uC\!W;.K	��v��0WN&o���Sri���&d�\ƚ�:�Se�4�k$��KO��*̻/m!�O;�R�yY�M@I\��j�aiV1�\Tܧ��s�����P͘lj�f%�-���$����"^cT��
�S
��� �B�j�^ʁ/:^`i��Hn?�t�M��BF���^���=�gFr�Qu3ʴf�W��4�Bd�J����$�����	ۀH՝�q��%������~��#(t����y(=�
��>��R�F��!�0{�A��a��R�:І�7jk�3d�'9Udp�8P�D�ĉhg��8%^��]�" �b���K��Mߝx<�C+?�K�#��}y�Q�B��.S�� FH�Z�+�3,�B�����R��[yn��4��iQ�b{�I�̐�&��)P��w��o (��$=UE�"��م�i�t��g;L����$�a��!K}:D�g*�|�nZ�'Aa����ͬ��(	�����V%��̍��%n��+��b�������u��oj~!%��#e������q���M���F�򳘥Ne�8�6Q�O��b�k=��>�:(b|��'T�Ѥ �4��lEd��D�c�0rx�ѽ��j6U����"�t%�"� ���.9��]�����?�^�F֍G�����<�[���=���,@6~�CrX&�f��{��m�����K�e�)�t�.r���kA��8��^q2{�"I.��q.,8y9^�w�bl������q�^����v	D���%�lȖXZ��!�N�w��ű�:�
�+�t���XGg/\cI�5��(���uE�k0��g� s,��%��W�6MY�_������Ҏ �=Ck�$Yd���^�ڿ��	��t����OQ_���<
+����1*�D(��G�0���}��Ԗ�،����\q���Oq�ov�9G"��h�m�aO��
W�R����^�Zo�٦1(�p�2Cyt�;�~>��7zcV]n@�_i>�	#�1�q#,�/]��I�kG1��.�l�3�������$F/t~�t uA�z9�x���zZ� �-|.rL��T�!3d�HF�j�ƹ~�v�ٳ�u��3�0���T����ߐT@�~(��p����l�5����x�9��<[f%e[a;���i1��Ҙ������[�R���w��'Dp�_򳺕�Q*l�Y��?>���Ri�eum��+���o���n��"#�/��`�Ty��r��j|��zADx����/�O��}�F�/���&B�w��~(`��vg�������,Q�e�	��&�oa��E���X���<ZX;�m��]Ppv�.�����g{����G���]���֤�8J�Ļ��C���M
L��:9J<QQA����g�0�yH�G9��ǆЭ�>A]")�g�B��Kj]��uc�����If��!{
���C��ӻ��k֓F+?�l��T��Q���^�."���� �P=��{_��|*/GSJ�������1a+��)&�L�J�!��},�½Q���7��s塎�`.����w���-�Ґ���g���B��*�&�jVc�~va�!�I�@uI�13��QwZ��u������9 ���A�z�S|&��>&�)j"�����R�Q'~K�"��*����p[�E�ߩj��>R�ig�o	>>�E&�nI; 3\���*�ieZ%�]�Ax:c`�Kzك>�OE��1�\ D�,U��a��{WyC��r2(T�B��g�E�?W��/�,�&��6�� ]���PX��?.������%��Q鵨�����3�#8f�K�	��@�e�
��]�����9�(W-)εzۯE��4�;�1>)*�J��<��|Xfs!:F�gݽ�5H6׏/}��\��ǎ��U`�,q��>�o��[����QKIN�x�y�؝��������YR�o�j!�](�+ X�&���1����kA����<�'7��_��E̪�
�}�2Ì7���DUS�����K�����&"�����0�#(.��z�Rv�Re��`-yG[�E��N���N ����m�@}U����ҪH�a�-T�`���.��,b�R��?��ʐ��8�z�B�m�q�Ie.L�Lv����NN���h/�V�}�>Ϻ��D�z2鋈�G=�v1���-��U�8�M*!���;��O�m�W��d9���4Jb^��<`ⁿŜ,��7�i����I�F��Bó�K]�-`ynz���=�����u�I�k�1d�Rhbq�_�P2�뛓"�~�׏޶T� O��J_�sTLa���@з�z�Jj_k���}6��(�5=Z�9�G�Rhy�?������Wek��Ǐy���G<>-X�WI�vf��ۄI%������cc$�XA����T��k�o�p�	J�z�U��G�pA����]s���Jc�ㄋ�GOU7��4w
Ȗ��d$�48�`B�y�~|��
%)�Z�ьɄ>|zc;<K8���.����Z9D���%ý;�m��S%��+D��Zz�L*�d��i�*Sϩ�Lt�ңP]�����G����祯���C�(݄����;L�
�ݴ8��@�AJ`R[m�n͔&q�4��IX��$�C��$� ��
̳�1�t�ȿ��e�u�c�V�(4-vσ��'����#�1�3p|O%����JZ��P��L1��4T�%�xJR�D���a�z��D�ݢ=pGN�?	=97���#��WL����kqu=��+�J5�UB���>������2|�D����� �'����x9E��P��{,�����%��L^��(�d9t��_��/���=���O"��5C���g-?y�a��s�E�����0d�*�)���Azxwq�j�KM��Z|��@�Uu>�Zm(�JK/��-~�N4��C��k���tGݪx1I�==�$��Ci�����	��_L��>�{�A�Y*b%K$���<��6��0'��4������M<-pt]'�P.�p������\�Hz=���ˌ*�TA�PrAT�\s�o�L��k�ozآ�?��.v�T4�������<��F
�?�E�>�nq�yl��X�zvԏ�V裠���..v	��~�	����H��r3<?L��0Kƾh�ma*C��r��#��?�0����`?[�K�u[Gl�$��
�%�>{AX�,�͐���ي�G��c�v�Á��0�az�hͥ┱�#�� �.�rP�2I0�?���@p�*<ПR�c��:Bb������-���sبx�~Ǽ�)Ό�?C�r��Z��'c탪)�M�Y�U�@h�6Ndhe5#8ׇ��صB�̹��O�3��Ru9��`A�7oR��X�,�%�kvbq�I/Q���lP؏
Ή�׍�ge2s�4�^�P��!G`�ӆiQ�	A^l]��!�O5䭋��B��l�8�&Uqj'���T;�/���TL�jGEs�S	�a����L�R1�7����ksep	V ���Բ��F��
76�m�	�k�UC��f��r�n������.2o��ħ��o�V����b��~r��A=Lz���Ĝ���*��>lO9����ZF�IT)B���s��R�Έ��3���St�g1�r��P���&�(�U��O�O6GL�"u*v�m��A����G0S9�o5r��3�2��Q��5?K�]k����w�-:m�=W�BB7���@X�����@l���MU�����AK�����h8B�B@�h�/4���7�\��U��:Y�����Q���oyط婦��&56U�1�:��n�Q�2#�#��]̃Ү��7�o�u֠����
vM�O���K�I/��Bcb%j$���<��z�g�l%��V�󵯜�2��'��w�i������*6o�t�\��#J̯2�`�j�=��¯�z�+��0�2*e�$���;�B�����X,`�>�C�n z�Tå�bQ�Dz%F�L϶����n��}�B�� (��Ƥ*�e�J��+������( �T<�]�@ڃ�*K�j�Zqa�>��j�|�	[\�,�YL���n�Z��J�L鵃��N��d���2d5�ρ�5����a%�G/�����p�����2vp���v�:�lR~6-�V :^sf�3A�&��x�2��C,G��x��0�uv�PЉnVN�Pl�Y�@���Y���v̥ns~9ťl��PTY*��Q��э���:]H���s��Bʺ�l	�0�����ltn��jOŲ
�<9�3�Y,��W�ɴlC(�P\O���ˎ�[�⨆��bA#��墪�}���#�O!Px�=jqX�]��.����B0#�2@�h�t�(g��;���<��f�I`X)���z�y�Ӈ���]�$v����'�Ct~��(�q(�ԕgD���:L�v׆�S�Ę�x�T�����3��6`�1�ȓh x��y�&0\�������!���E���`l�i�B���p 
����yP�a��
j��4���E<�
2GIw�>�f-� T�\����rW7|�VĂ�×��W�mdv5�e@	�d��e#+΅:%��R)��!<�.�U���K�60�u���c�"DL���(pI&����]Y�;ó�R�ٟ�y+�]��{��,��)i��R
��Z�*XǄ@��8�c(g�@�8W p���]�nƭA�O��g��B�,oO��������|�Grţ)�$2���Mmk�-fCu{CU	�J��}�����nu]PV��Ϊ/㭐n��큣@��0X	_�4���b�%��8��ȓ�s���t6v*K�Z� V�>��n^z� lLޔ���&B�ں�F���1�o�&�.:��58��w��ϖ�7���0��R̽WiH���^5��n�A���,4�-<G��w�1�80XX�ϲ�!���`�ߪ�8|�y��Y�]Sxݘ�Y���ˉ]���$�E10�����fu��ȡ�W ��Ф�9�TM�zݿ
\�����?��Q	��2D�=�ϋ9}f%j�嗏��̡ר�Ӟ�F�k���_���򘰕!����N�������@Iqù!�w���r��XS�Mև�#3\�{6� ��O/�����c�4E,��؀H�j����]ev)��"�4���R~'{b�%��Qj{qi��Aw���������yТ�F��r @$1~ʊ^�xSv6��o�f�f�R�x�;:�}r�\C�⿋Y��{�2�(Eg���T�I�e��O�d�}9si���'�%��d�����*v�����q�(�A��P��gA�ϗ���juJ��C��
*���<֮p�=q����$�S��=�%�N��"����S��y����B��Bx�)S-"���7�J�GN�=n}UO���
j�X8#�%3�ߒ�*�*��S����ߔ���#4�-|�<��i�{�PƎ�K�ˑ����N,�x�$񧓠o*n:gʸΉ�N�n,� �dڄ�P;H�/��y��5�QP�,ʱ|��كV�,�,���3�`�y�[p�hpf�y�g�D��d�#���'��T�6L�]���d� �/ ��qpq ���h��dpIn޻ݟy�d�u��@�|�;&�
�Ey���_B{T;ZB��T�f8�)~Rqv�vn�����Z��Kg�b����k�:��2^�qc{Z�:+A���{���>���t%����(q� V�,��F3Y��no�uF�WL�Ǩ��4�<���p�E3�ta2��	��$W#����ŊG��$�Cr��bXsu���S i�[�|�+�`�:��% H%��5�_�������`�y�OX��n�g�
�|��ba��,� £�7���Nxɮ
@<"g�P _��PΡ��]����fwI���K�c�V�ݽ�������N��F6<�-�4��+S�)1��o���v	z�,N%�����#oD��_���;�
��%!A��\,��΃�H'B����3�^u:|VbdK|�K5�u��s��� �Xa��驠|-�R�EVg�0��_��+�f�{	[\�՜������{����$[x��İ���N}���Nv$EO�ԟ@��u�K�{ѣ@�w�����v�{�AF��
���vV�w����qW5ķ����Q��SB��<�.32����:�¢���c���Z0>�Z����O���x�u�@�����y�S�tmK\N(�Xw(�:��k�j���⧁c� |��̘�|2��_k1	�mC a���£�r/-]M��6	L��ߊ.Vsc s[쥲��w�%�݊�c5�7��F���0�U^�2���l3���>�H�=���ٚ�=v�|kB�㇟�ALS���_ll#爾̙��L��?yXQ&M��[
�7yL �7k���TWHcDE��l�[��5>uɳ/7�D�2Kr���{-��/�����R���<5>s;�7S!����q�)%�f�� ����@l�~����-J�"ZޗD�*��豬p�0~HZ��`�aLW���ko�J��Bfs��v+���!��hw:��:.~��X��74+��+�	Y�8)�5�O�c�t�?�|��]n�-�R(;\�#[�\3�Ξ����θ�랐��9,�XH�]C��4�����3�PYP��n0�3���Y�z,����Ȁ������	jO�{D$G�}�o�@������$��c�G��B�.s�@�R5���	Yƛ�r�vU�I�50���{ #D��A�e��j�e�Ϟ�'�/ǯ���a!MP�c�Z�jF�Ī�ݷ�#����~k;�o�&qm�(�GY�Ȉ�*:�G<�=����\ӳ�D 7u�2����c9��d prW�l�Ɛ�E�b��G�x���ynhu����-�@���s��p�㫇%~2��H��_�(ű��"2��Pa�S�tI�-s�QU�O�&�pE&��BkmS��hV@ �U�.L��!�א<�.�$z-��G��P�!�&5��& �S�� I-�z� ���Q�8��_���sE�nT���=����Mba�UT��.�T�1��x���2�V�������YP��s��PE�:�Ŗ��(�ċ�w�դZ���l`�W����#�
�\%%3J u��hJ<�mu�U�m9��T��^��k��e%6&��k]u&TҚ�����]Ra©{�7�0���t:iG��uR��q}^����+����YI�e!RPRˡ���<���{��f�uX���ԃ.��|��&�O�;%E-lUđ��m��4j�"�����X�h�u���0R���E���R�\]�]Iv��3�Y~R.���7��.<ܱQ�C���cⶑ"a�lΜ�/��ch�]��ņ�ʷ���<G%��Q){.�ޯ^��\��'����N�m	R���m��n�������q��Q^�۳Z���/�c${}����|Sg��K�1�ȸ�U����
�RVV�3�;]iG��������X��\��B}���c;���v�����$���{��z�]�M����6��#[��qO{��~l���ϙs�̻?S����I�eo��	��K�����E9c��.u��:��;/�P�� �3�ܧ��Hp�~��G7Ԣ�ba{K����s`���hxB�G�&>�)BA�����0B��m
`�R����hS��:�ґ5���xR^F����*?���=�I�ɉ����Y�lxb-eʦ��U�j�p�L��5���==���J�.�=�Û0@��]��=��de:k����Efyf�y���wM�5%o<�Й�/�2G/�V2��U<o��Ѝ3P�j�۹w8if��FD�al�8C�طy���1k�H�G�Phc[ώ�G�*��Ȁ���|娐�����1�T��c�dLTV��ed�x�!�B7ǩ@��	���^�~lU�΄���Z�'��C�p�6�L�*D���;��@���9�`T������lm&8r:y�~��t��~L�|�CĆ����Aͮ��d P���_j���k��ݗk$�\�͔|G<�r̷���";���:~���V&�N��D�� D��B����)f����nQk�ͼA���}IUU�R6��9��o��4焹2УW"K�h6���E?�h�������t2P}����O�to^��a�yO���Gq#�*`Y��R�Iگ�-�9�2E��ϧ=�5mJ�N-zכ�0��_R�g��ۭ��%��4#��`Y�͛K��ƌmA�o���=���\y]�UKi�-R�2_J���U�7nr����ü�D��0R��] _�bgc(�er���f���A���66.{����
ɆǢMGm���`b�bY��,W�hz���	5��g��K#��1�����g��/�r��9c�K|Y"�2Y��m��>�,;������0�JL�Kg+
z����eQ!�ow�%᰻\[\��蠃2��5�'�phbM���}oNn��!�&"�Č�E��<j� �'5V�+.��:#����˥!C4��R��}x�&��~�&�x�MaiV7V�ye|�_	�O�*��W� ��ܞ��<dp�0�}���]3W�牷׽�V����w�t�m9UG���^�&�/���w�D��=lʲ\��s��U'EY�o����.���\���sX�8=����\GD��h%+��c�J�P��]dR8*�߳(�(Q�܎3��������Y��_fp�����;2�Y3����1��y�C�߲�����f�l��@0�':r��������L�V�� �y�|�R�Fy�˝o�C����F�.^+�ȴ����1a��^��ώ��0	W�����V`|�e3�&gWf���LT$�_ 2|�	���A��t% 	����nW��C	`�7ґ�X��Փc�|tф�#�����җoe��_r�P�jx[Þf�@�8��R�G4�]���F��;��!�]���j��4���^eX`<�K0���}�^�!����40�RX�n�x�R�a
 ���\LG�fv���e���ɀUHә#�LEF!����o��U��<J<y43�~Pj�Gf���9NU���k�j��w��?RޛM�K䕺K#�������P�;���Q��A�ߪ��G���q��5I�!�"�a7|wi���"��R��XRu=�@��|/?�?'�����ɛϴ�`>�9���=�h�Sw�`�A��a��ߜ{�o�2�>��&���
��w��A�k��~D�b2�d��;]D��Zh4_�+��|
 [���w������Wn�ɪ���tS	lO�5�����r�?�hf#�5�O���'�?��Hc��cJ���JO(�I��-���e����B�>��*
�|S�e���z@rv�c8�.�~�L5ss15D��*T7:�耓������"p�T�$�]$iN�Z�$��]�m�[�u|Ѹ��� �C���H`d�g�0�w���b G>	�*kr��rdİ!���Oň��#j�4�KQ���D�*{�3��-�l�՜�D=�p�
I��e�X]�|�2�ᠦ$��8d�to�)�T��w�]�D����;��6Ҏ����fo�ƛ5F���K���0�W��Е4��:�!}P����*��(Z��E���~*rZ۔�K� �ǝ�ߵоhͤ��R�� ��g�����Qܵ!̞� e�u�X �!�}����fA�����U"�&0���{��$�g�9]>G��q���K�Be��qF�z<j�g�xR|��kT��3����#��4ŗ1v�zGr$,+�2F�-�!݄i�� �O[�U��K��oX�O�6�1�B�>�,e
�C�M>y�'�	v�E�_�m�oJz��1�W�-gm��L�������j��MV���5��~���-e��a�E�w�.&�s-�]T+���t�zhE�A��2'P�\O�.�^��E�6D/?f״���|���L�1|�ɬ�1s�mb2>��H��o�*��o��f&*H:��y�O�E*H�[�ll1�9�O��&eZ�!�zCBXZ��Xύn�1������^EJn�\:�K���v:l;'��oi�2gA_��au����.m_�l���Pq�:i������j�&�  *���l�u���ys���+]:��~[�q^(����j�E��Rʽ!�A��H��3�����U��s�'�b���/��]X�j��i��FW *��"��I�Q#L_p.�pZK�w2Oɡ��W��SM��%���z������s1���#遇���}�+��jL17s�d�{� �F��Γɿ]p�y�Ό�D�Z]�r�F����K�K���P>/lf��9J/�h�W�#~g��������_��,��,��? ���[���{ΧnV=i�S�,�����u�R�5�R�/Qr�0ϓ=��[�Ԑ��M��IKY+{;��/�9��؏H�@x�ly���n��<��������$"i@E����Xia��Yt���G�t�y��D�	P�Z�E>F�TYY��s�5��:�����?$:t�Oξ�O��K�1{�X2�ļ^����t���9�Л�V��>�̜ڭ�8����K\m�H���8N��`]:���=8hUzlg��$��)��wB�P׏Fv���`��x�N89� q�;�!�h�;�l��u+��>�'��`�6�9o��
����N�E)ν�T��3gS��U/���+8x
�@��Ӥ�cc���6l��8�� ݶ0@L�7��A�E�`������&k�w� ��TnBS����]V��d����_	�;��L��X�NV�SgRG������S|
	�g�?��w�`�|dX�>����	qb����3o,B�C~�������	�͔ ��kaYm��V��xY�ѽ���������*��S��$�Rg�J�����tm��o�Ύ
�Η�e�6F�"vd�J��N�Z��i�L�,�Ptxr�)���ƹ�J�`��÷y�GS�aY�ꩉu�F3�G�4��a;H���J���/��9{Վ�dBڜ��,-����ɭ���OM髆i~qc$4(=��zkĵ�|m����+�)���.��$*s����]#���	+ڷ�6�j�.ч|K�[�х����q<+Bm�\��RZ_Jk��a�I�]�*{��іK:�;�
{�i���P�_i�;��^���2"�v7���9�R$I���tc��[��7��s6��(Jj�`k�/(WlC~Y��[��Y[��z㌏��-��Я����A׶A��-ڝE	������d�r�%K
f��#	�J��m)�G�2��"��am��X��+�	>a�w���^���ͯNU��\W�"�޻���)l�b䋭�LvTƹ̀�u��u�� ��~�wb�Yє��naS#����{�oH��9�(���J��g�<8JmF�uŦ�7��j�$eH����|~�c]{=��N�� �{.6��~M�M,�����V�[�
����8�����Z1$d��B�l��π���q��� ?FOB{$�,�oӛ\���Sd^J��.�t���5G�$����*�/�j1��R��ē�a���\T����R���F6��#�᧲n���DmM�)"��l�YX�� �m��m�a*ۏ���n[Pn�9���{��4��O~q�R+ �A��k�ϯ�h�{�x�?jqE>oK�¼���y`ͩ��d��cw>��_&�(���[�n�.H���	�	p�^�а`\���BR�7��a|��4���鞟d���<3L�x�[i?@��-��2a����=jԪ�Mo2b�֟�.�h�(O����2VQ�� &Һ�鴪�������w���o{G�8��O7F>�����r�ɲoQ�K��cf��82	�TֵH���I�Ls�����)u���q�ŧ/R�(Z���&��J��Y|�X�F@�6�kf��p��:��x_)d���N�� ̫�Bm�5�'����-�{���4�mE W�B��u�ޚU�W�_8��A�z׷i�]HA�$IUM�{��C��T}�����
�H�w/�cj-��Z@nλ��.w�I[U?�jA��E�=X[�kY�5}�O�ZSuB�#�Uh{�{;�qx�I�
4�ScD����ɻ%��'`�J�P���V����3��fN�L��Uy+���ޥ�����U�c��&�,^YH[�L����p�������S������vZ����f3�?.�����t� 9[�M�T��M� Ⱦ�7�&u�d�L{m+�L~�,֖k�lJp��s���Rы�.�&+Q���G�Tm��0�֫��n�q������Uy��_H�s��t��q|�՘́�(s�+�̬cۭ	^���"���L�2qݼң��*���:�LE�� ��B%2VR����(Z��,�!k|g	㒮-3�E�hRXV��{B�V��r�K���x,�^���@m{��-�ǵ�\U�yu��LÑ%��k����|�f��my���ҢGco�bs=��|1����^G;	ǥI��|�����v+�l� ��8��F`jF�;9$A��Kg�}5#m����to�! �kN��b�c`�UnUK@�ˎ&�8�˺�n^M���|?�n�+լ|�P2�t��J� O����������iFc��HĻ��qY.���,P[>��K숙N��{b�S�͚�n�RQi����S+Q�p>b����g�Rp�"���?��0 ���1.��f�2Ч�F���R>���c���X3��_ޢ3��e�lE�7��E}��7Jr����\~q�ןN9����*L4�������қ�����b�q��Bf7Xi��E�<����f0�ďL��'�����;�ю�k���K?���JqVM��*�ÊH/�f��]~B�/�������3�K�L��m��̵Y7]��_�y�Mj¸�HƐi��^�+����;%S�� ��.B����P��-��k^�&�	+#�T�
����O9;�6w'̈*�V�@��C��w�2��ռz�h�	a̬f���s�(��ex\6�奈��ԩ�t���p����!ބ���i��{M���9-�K�1�n�"K����~	����~�t�Dխ�3c|�+�1�.P�(�֟��"�a����d��ŝ��lg�e�6(�]Q��ķqh�W[ʄ�=B�WY
�%��`Kx� [���uK��^u7T�w9�(�R8KxN��7xutz���T�� �R�n�,��,s��U9q7����:��L3n���v�� �����`��܅rt�C����<���1��Bo��W�C��[FT�?2�J�rL�[Z�pcA�����禬�4�G��^rMX^³Q�<b�=>`�5�S
y��mL`�Ǔ)e�S����d���	S��RWA��|�:�'VU�V"A��¥٫�1oL�ò�6�㘬Y�z%�̣_)����l:j�~`�q�+o�T��"�6�{,Y<�;rF�T�`W���0���9�?O���z4��y������z��C`#=��]7�L̐=�P�Яm�.B@�G����Zn-]�T�:
N�TC
��)�x�x3[^��z�炎�[���hˉf>7H��"����!�~*�r��([+5��1MX�Qo�.��|N$f�|6����������{CĦF&J=����n3�ϸ4F;�z�#ԭ+^���+��8SX��[�"fC�"s��}�@o��~��������DZX �$�r$���B.�WR�Ϯ�S�0(��&a�����P�4;��1ĝ�&0}(�uL$���l�ϯ���6�<�1�R(��W�#���E�*d��z�q�n��w��r|���U�݌��-v;��b+�:�"�sÐi3���&��;�B�7���y��\�ω�_e��m� ���k�Y
Q{�+r'-���6�d�Mm?�JE�h �w Zx�Uy88�܋�38����O��#>��슀/֊�����h�&z��9���sΌN�����<?�`ǵ���:2q>w�����Y)�覷�Gm��M&��7h�4�;�K��ʏ���BHҜ��踒	�<'@��ځ��$�E��&�3υ�rH����΢[�o�PR]���?;��r��n�B���B�-y��$r4�����ft�[qc9;�b�������������@��g0�Ԓ�m�-��H&������*`&wU1�
�X�I28����߀��M��{nH�,:��gD��;_PLOF��|W�i^�.���_�r�ٽZQ��+󧺅B�����G��=1b$)�^ҾǶ'l �ͤ0�U�����}ܸ#��U)���|�E��.�ؔ'd�Z	x��v!����6�7�~�@թ��o;�+YD�Cг��h�{߷i`!�h	Dt&�M�!��_���뒷�B4PY"ʹso�"{k� [�F�/���p���]��M�g�~.�H�������Ƣ6m" '��V��f����5"���XI馆1����KǺ~��'��|(�Dyz�/��G��$*>��$��L7��+���W��e�S{v'O>�j������r�E�{�״�YP��<.�I�T
A=X�h�L�8�B5=g�g��X<��9H����So�BxOWp��fD��b�Gjs��V�T���6p}dֆ��J�Y�$r_\k��v,�,�k�v9�+39�b�wc�r@ʏ��3 ;�X����.!����c<݀yA��8$�u���N!7�D�B�R���y؄�nOc�(�񕇒-����=���}�F���C�FS�����Ŀ�v��<���
��)��DdĤ]%�Ʌ�t�7eZcH����L�t���Te[�߈�d3@ȓ#Zك�Y�S�܋_��ó����j��ҽ�J�Ѡu4�ʪ��'�m�NSI��Йe�ϯ�Qsy.s�;��+�F��p���ԗ|�X� )��'�d6V�49�M�	w! �kM:!�G͉>��NR��hä�)i��5,������/�RU樉�^Xz�AǹJ��)��;GZtt|
=��o�_��/#x�A�� 7<t��pB�������Y�*�6��RC�$ X}�F�oZ>���}���C�1(��Cs�WV�h&q�l�S�L]tM�În�:�3�X�у?,ԵV)*�}��q6k�obA`"s~9�i7� a��ss�ӯ~>�����%�����e`��և����/kI��n���s��qc.-��
*-��]��;���)� Y���	zxs"d1F�����<S�n5��Gn�cKdn���}[�^X��Ȣ��Zr�ʘ���GA@�`(D�c��ݦd���^:/���u#`�{�ȻF�w%	=^m��ɔi� f�n}�t��D�oꃫg�S���^���=[�C�x������&�Q��De���Q��!C7.aQL0��ظL	}�0���Ҿ��X�Rq��d���f�s�����@z�X���a�^�ǭ�,�9ݎ�6�<K8��b�;~v?�&�����2R�[)��/'����_-�;�JF�C���c�W.��F�8�q�J�E�녽�(oE�Κ�SVly��e���� ʝ����+��Hٍ��w��Z �l�(�@�)��ixXw�l���"�N����S������`��7��W�,�mƩj;���>�(wx�0��]̍׼Iώc���>�
��4��òӐ%eq�r� �H���p�63�umVRG)�������A�B<�^ä+�ѐ���|��8�PH���B$��P[ �Q��Uތ�jgoi�sʉ2S�E\@xN�"$!캥��S��q���������4���'���y�j���$��=���*���/S�%�� 5?b�[�̭84B곶�1�����:Q����*}yd�l����-�����z�B��V��1u@i� GP̃BVOsG�������a���� ������O�����ٙ�8xO�h�@��-i-Ѽ�4����fQv����#�Z���5;f$���vt/S��?M�����Z�(�G̅x��Z���v�L�	�6����t�#@���0���#|(��f��.\j����Oz2��(i��u�VB��A�ai��V;r�\�cLP��8�����\�x�m}��z0>>�C4�ifҔ��zH��	�'�\������liPq?�ӳ���s_���Zp��⌉���G�bG)�k�$W���"�-���X��������r�݈yh?��+U�Ґw�Ks"��F��H�ccy�4)(<�,c��Őp���H���Ɗi���;�a�ځ�e��Vl]↭7)D����k�o65,F���UbPNA��xR[p3�̳��7�#����T�^;ȯ��Y�¬��Um�o�c�_�k-�@�91�e����w�P�C�l$�$#oEy�T���ʗ����g')V+�\WS*��ޕ9� �*�:�~�wϱ�;����ȱ� �
����pB6צe��������򺏷YQO.z�Lk4��W��5P}�}��V�RN��4�Tu���T�H���>�C�զ�����(9`|�x8H���:0Z��S�:�������[�[0�%�%���bIn�F�e���zk��-s۽1&�k%�1b0���)]�P)X(�r &�"a1�1���A7�W(+��L���*r������[�����hM��Ϛ�iz��iC��4/��D)�<]���	I�@+��Zg�餁����y�����m*O��^�g`'�xd�_���'`�/�JՊ��?�P_�8Y%Zۀi-=o\���?b����8k�GԽUfCӹEbD�H�ku2 ��qF8C��}�AF�_p��� V��h�}K~��ok++�<$�	=B+��ɽ���*6"N���́��S�����-�����pL�M���= ��Sa?�C{Zw�!�"*$�9YjO�>�s��p���o4l̑�b��5L�Ci�;@��N��@�X5�=�1��YM�م�k�w���eY�Ǘ��Uo�<��r��,9_t�k%pCW>��Y�G�ejU�@@�}�/��X������
5 T_�J�?mK��$�!%�l���!�
���тC
˭œ�@\d�;,'���/��Eٖ���J1,b9�p��e*(�������5��U�z�w� �n��ź�wk]�E�1��A����]��&CϿ��e�Us�xԱ�j��%mu���p�,1Bn<�y�&��O�w���C<��.�ٗl?j8>���?�t�����
7�҃�/'7�%���d�O�Q2��
�rh��B%�r��s7^�`��f�!-�T׿�h	�3[�O����m�<��(���8C�'5>���,���޴�w��!�lj��J@s�� �D����G������L��Q�}��Ϡ,��?;�Q���!�w#?���+�T-��u;"<��	�|��0�Јf^C�R��U�W�E}q#�rP}�aE?*��z�P�f�/^�����-�U�
v�fߜ���IXGk�!~�"h���~*Z+N�Z�܍Sd�dKM@��yM��1�z�2�spK9;��{��h�A���rCL�l-!3�Nh�(	;w�u��mAY=��D��I��Wb̂��}�9D��vp�(�*�pz���'ӹ3�(�F?"��/)�A�����T����s�>,Kf�b6��{�|��ƻ�:3��6!���a��,�Z��̟ȓo{Rj}��R.<�F�NZ��Mr<K�6�G����q�'�*b5��O6�V��5�h����6��?4IM�i�F�i��&��&i�H�ʾ�������}���"��H6��0��cSNH�U.})/N($���7��ֹ��kЫ��L,����sL��snpzg��
���#!�}%x>�A\����n�{~w���a�ϵ ��̎4�g�� =�����=��� ��T[��IU����{>~)���^�%�	�P�ȑ �m�^��B��i�T�_
綰�OGJ�_��"��H)�V#Bm�&1��;���3ä�G��6b*���
+����`-�3�F~*Nԩ��*C��w�a|�a�%��(�zn���X0�16����:����.���t������V��pމϦ*-H
�4#�:�Q-�]G7aB�(/�_O�!$��DD���_ �b�Q`mg[�kn�F����ܶ.bO����D>�'��?��ӱO�����r]��y��:�땚���?����$�}H;�t:��bw� �N�fB"jm�h�X����X���;6����<>�Rmٟ��yѝ�@��J!���/�9���Y�u�dh��� ��Z=8���B)�_�w�~X�?!�O��i���z5�(2g3}կ&�*H��E�� Y+�5��Z_PE#p���0=c�|���ϢV13�G�H� �O~[���D���J҃ $�H�ЈTE�D�]��k�k��[HA�ȇb	ֲ� P��oO�2�.�L
|�1�(��ڔ�jjL�Jt�Q.65J��;��H9�#!+d֕L�I��}�KC3Ƒ_<{�^��f�SAt�<�o_N��e^��u�rD��O�{+���=��p%��άņ,�Vr?!.>\���3�������1jvR�j^��ߤAK�Oa�1��UJ�䤾f�1�K��Ds�2v9hgT���Ί���R�|���s��Y'�OĻ6'�%�����#�}Y�Q�
փ��$�b�7e6�"8��$�ۅ}���{����Z��*�îpz��&���F{����$�|SB��?ɩŭ��������5�/6�@��1Ǟ��"�r����1���>#Ćh��V&�Z徧V>;��DWL/Q�w@�'��~���椺5�Y7L��ۘx醥C�β��ʂ����#`�nᒇ�h'5v�J͛�Hs��P3������G�p�M��Z��riii~1�dhu���S�Bv���]��Y6p'l�����ҩQ��b�썎+`8d��09�P�L3�I[��5c���̠�q�a6!�kaB��,��3S%�_'���+r4R�;��ԋ�|D��R�O& A(�kv�BZ�����*f�5;;�w�[�UA�˿P4)⹈(VlH�!"˕	���ޢ���Y|T C��bJ�m����Hڸ�(*e�G�Aw̉�!��m���>�l�W��2ZaS�l���14���m�t�+��;o�����ɥ^š�A�g!8��M!,��摀+�`y�'BA^��TͿ����������N��Z&�__K��~�����5���ǵ���è?3�;����;�<Y�W���co�(��TN�)v��8��ֲ1ؾwWz��#/m>]`N�����^�����e�����+�aA�厼�f<{�\�'��7n���4��]���.����Df��$��h�,���X�-Q}דP�V�yp �@��̃9����蓳CWhp�������[lf�שzr���E/c�C�p�n�0�}��@�d��d�hzFM���?�l3H %ݐp�`��<J��`ɋ�6R�����H4�v��q�b�+������)P04G�� P� ��O׽�Wkյ���G}��a�j�����J8�(ww��)�Wkjy1c���[����Dr�\��������Y��Gg��ufI�R'�?&/�}�4��d�yh�w�f�/+�b�ɞ+%)��ё�nI�8VM�
B��� ��j�@�w�H۹F�����ұHR�q��Zl=�ڏ�F�#�v�7�qX�~m��:�Me}�������),�ڪ�g�W�'��x���. ���������bf����?D����2j?<�� �\m�9��;� �E�ҏ<E� v�̴+�
k����E:/r��=m��YSt�1ZVQ�h�)r0-]����9�~���ۍ�n�п{�����xI�V�a�?$i�]U���~���?� :��ɂ[�O�d��)�#�P�t^}�Q�����J��I+rE}�{���;���x�"��J�H����	�S��#���[����d���m�dBi�|I��0��~t��~qn�w�u�Y��bM1,�S��`��v��9!UR�mB�����ʐ�eGcTB֭v!� ���A�plb����G��;��a5�^1�]��� �[J��Amk�Ջ�?��5���S��p�-Y�Ϝ�\���S�6�%1(�ߺ��
v�w�f�!�E�&4Rd�*�lLǨ��G�#2�sC/dgY�
K���Z��]��!��O�P���yrL��[�½uU�_�d\o���(�4��k�%�pf�����\�\�C��([�*>B�;���O��5�6������c��a	;���D	:{K�Si��0�C�W��_,V��| ��D�.C������Xv}�����hN��˾�D�K��	�'�"��xX�2�v^Uk~�����EG�4a�����m�RHG[�/פ**������c�^�g�ƀ��Bf�25��;�8��b�#������R(q�U�z�G�����e�4�\��֌;6Ϛ��n���H��,�����Q�躛�⼖{X�񷅠��Þb@W�"��C;!�g(7Jp�P���)槨��n�����&��I��Z����Xd��}���/��w|��u"�CAB��ſV��O�#N1�����s�rT>���{Q��*��`\`���!�	�+u���q��6�=��ԝ�t�	)u������DF0�
�w��k�t^y`��?)�>�R�k,�f���Z����¹g���[=\�P�:sO�^T�x2�6�c��P��[dD̺�F˃���݆v(�&j�F9�'�Y�⿪�q��%�wh�	�;�[0!��X�8J3�"�-o}�ܧW�:O�-l�.��mt��>S�����-�����ż���Fwk暑�i9k��PE=ޘ6�pL�Ӭ�ۜ�5v�M������m��O���ⒻNX�R��{Q�J�#gt�ӌ 6=�oH�ȥ���+L�Z����إ=Ħ	���`���|�m����ᨳ7<�/��!����h���_�1�X��a�i�ߗ���v# �����A��X��{ ��>޺뽋��	�g��m=*q[�6p�KXẢ����]5��)KK'<lݾX�WxНM0$1:�Q��.���~}tG��Q��x����HAb?D@��E��-�u����Ea�Ot@��r�S8M���t�sVM�8�������^OE91�gd��98�[݋I�fG�q��/?�W�gPiH�? ��l����jb|n?s+�q�~s1T	���.NGz�}������@A(�@ڣ�Ͳ���(���ud#c@��?ˁUow�J�ֿP�&���?�o:5V��+��#��$˭�7H�5ӫD�Eҁ 55�9�m0��|L��`��`���$>0����|��K+�T��6�kJ9���wF�P��ɕ��Vk�����m�2��Q���qX��5��"c���_:�X��(� ѫp*�z�GCr`����wU�{��<u��C�������d��¦����J�Ǖ��
*��[B���&��ŝ�Ɉ��E.,���F��������3iQ�1����w����E.-��zJvJC�0s�,o*��~��,���?���[���.y!O�6�F��K/>�641��7L:���82���-)��>Y��O��hJu�5��E�?�_	���"����V��h��P�p�?����	����p�w���<m�ʇE���]�	�X��Cypo9�ƴ�@:1PeE@?��㺜sN�k�3S�S@/v�P_r	-Nf,H��� �NJ�+o=P���}r|xB�/z��oV���� @I�zq���'�U�
k�R�ji(�#2�� tZM_��y���G>�yg6QD�)_Q�G ��"��{�/l�4��7�"��xKH���S@�Ȇ�w�rH>3h�}�Ag{�3s�yE��Qc����uF����Wc���xW�l��(G�w�؊�񴹵�P(J���`�$�H��
}z=�����،�o�5�ȥ��!��P޻F�#���oo�R� l�w6��W%�~�A+|E����.ؚ[�קC��'��K�s\���U�?��l�5����q�5�O�W��WlЩ�R�ʜ�Z��]b�|�x��Y*�w'�����D_Y�ֻ,�����t����y� E��0�?>]�"�a����_&���ꚶH�%
�i��'q����p�W�t?�
i�I ��6-��v�ѕ���E�hOEA�8ץ��8��0�7������%���Y�S����X4:4(s�q��v|��m�=}���V���o�{h�c�a3��z
����aCP�O>���Ĝ�U6�@�Cu���~*2�	���{�����| h����h��߷�r���T�ޔ��Sa+Ń��(^9��X������EmH����Or��D�$:�:�E.�e��9����5��ݪ�`��[��������
����&���P�(��-).�����E�7faq��7�l�����p��b'�"`������b@%?�YUS���It`�{ bo^���U�m�F�V������p�O�d'Q@�'�7ұBY!�Jb�#[�����t,�r��޵\>}������P�*6��%L6���5��Y�-�fi�_7o;��Z6���=Ʒ�и�Gˋ�y��t��	y[��e�a^E�s�U~y$"v�,x36^vL%�7-�$�؟����,�Aaz@Y7�>t>n���d��;0�v��e��p��Vo�X\��exMU�d=	ۧ��h�59	������j�N4�[7��
i�K$4'P-V�"��_�ezu������1����� 6��:���/�.��N`X�u��
HS���`/���s�ya�������Ea_k�5"R5zU��e�W����58l{�|�2<E��՗C���e:]�򮼅=�Mg@�H,�P��O�2��Vj@DwWW��M,��,ކk��8:�;k����\@Krn(�W��}���p��d���lB�Ž�p��m7ˊ��z )��D�dJ^5�����r(��Mk%�eB��]��p���|�hj����=�Ê�;�R6�|��&]�f�w����\���(R��u�8vճ����,t� mm����  ��t�*Pt3��ԴQC`�*1�Ń\�#mcя���t�`�bA��\�_K&[�X�_�+f�,0����ʛ;��x@��"2�cɮ�R��+x]�$R-S��'Z�9����&n��U�ǡ ��ĳ5�i�n���	������ܠ��$�� R�"�#Ԥc� W�`�]7�W�O00ms�N�Չ�]�����˱��!r��wi���� ������,fi������i�0��MH-k���=
=���۶Q3Q�Or�U��kZ�Ho*#�6���h�E�]i��N�BO:E�2#$�]	�s����QB�yN�'�K�&\o���?��|�x��U���K�R��me��ڶ��L�``P����HL�Յ�T��Ms�3��i�jk��7j��/�k��i�pW&�cވ	����`�=��=��i����+�V?"#��c	ڍ���s�`锕gh�y��"��y h��	"�89�R]���s�[s�Ӥ���Q��6���$u(�� J^��jaP������]�p�!֨��d$Q�Pͷ [��/z�6#Ã��{�*�%���^�^97��ڌ!�B�ږ���I0�;Z�����B�ߨ�؛�5�h�ƨh�=ѭ/4���h�H(Ji��N$��]"���<�G�'�-�����ǋ����[f�?�Y�d�/�f�X���3h�p�����(b8c.�	[����6�6��%���4J�9�N�`slț�*�#t�V����`v����=�̦�t�*h)y����4d@�0m.�����-��%G�1o�)H��=h��l�վ$�@s�*��,�
�Zq�F\�&ǭ�[�//�V�`E��6ڵvj��N����� �#�y��X%Y;��l�J�B7�{�X�f�+�@�Y�4��Bw�-V�-Te�fh_�d�\�d͎hN���*3
s�hB���g�X�/�/��&'<Z�[)��賌��K��0� oh~�y��B�o�=�,�`���h7<��#W:m|�o85���#�'E�nv������qW�+���?�c|	�z����ٍ�g�7/w�~�ڲ�a~GNպ?_��
����En
WF����C� ���ɞ���b�D<K�
���� �kǭ�$�%�n:~^� A�MF/秙�4LAy�#gՠ�{T�1��~�0�ԗox@@��J�%��Gp�� ���ooI�(��̛�~ֹ;��PH)r^?��yZp��,��pK�������ݧ@����������5",��G-Ǡ�ox����iQ ��O�rVdb񘲸�2�n���4�ި#���/ >�`;	��:�ԃe�,�c��������V0��5��X#
l��}��S�T>+�J��_�fڼ�OP�?����1?σӖ��?A=~��,�k�vǷ"�^SQ��_e����&��`�r�?Qy�|��X�􊺛&J1Y�`��1PǮ6a���b�r}L���"F.�'��eȀ���S����"uы���&m���ۢ���l�;�ġ5��8�Y�]4h�/����u&�卄�o���e�I$>�1��`u�|I�u�O���saJ>�W��f��T��WQ�=�?j�o�O8�%j�l�t@�Mp��e�H�^���jq���ڕ�y׷��.���0���ص��zܑ�!�o.�y��X��Y!��S�����h���x[�Fp�X�ތ����Z�&� ��-7���67@}���i���Q����E`I��ATzҴ@U� O������KB�v�B+�k��}?�k��{�#.�U��A0�4K{꧞e^�g[�b�N�uIP��cȅ\Ǳ��D��w_[[�%k��m�	��Kq4���^&�KޫhnGǿs4m��c�V�;�3˸�s����A�4��n@B�-�̓��GP\@>����AQk�N F��ޑպA���JԖ:R�3"a0y�����.0J΋��ˉ�������zQM%�@LgO��0�-���`��pb��{[m��驵y�jR�0��Mh=���>����phkL���U'A�wc����M�ە^��%{����O��d�낍����q�������.b���,7ǟHC�X�A�)	�-T���.S�S�}a�t�|����(������6�[~F����M�/���ϱN����G~|1�$�٫@w�g����r/��s�
�'d�9��=�D^~\�VU��#	��h0ҕL+���\G�Y�`ZU�-���qa�{d�mF��^��0�^
&/Q�C6k`���_Bg���nK��~���+_lJ�L�%�_$��Xɠ�?	� �L�����T���Z�-�H,G�h�W:��n�-m�� ]7:7}D}�xPlQ~�l����� �K��b�g�sF���ܔ���j�t	����ڻn��:Vּ&���~�_� �{�QKf�D�0����ֵ*���u���=<�E�i}/�G�:����v]}�d*�m���:�L5�;�;�5#><)Ր�i�#����lN���G�[+f���v��P)�aC+�9:������2��T����\^�ީg��f��ی�Cш�n�â�h�ڶ�Y�L������#�{��*�I�B�'���P��7���Q����M:��L����7�F?e�Z.���1Mք�!��Tl�{:��y���9�bT�?ėk~���!txCi��(Odz\��-��2!�uhdY Aʉ
��>���,�ob%q@G��ۭ�׉θ�-`Č��R1�I����^����~��A"��x��e�v�H����Mehܲ�x��ҵ��d�l��>����x8�E���[��ۘ<�t@���I��H��O�ɻ��v[(="��n�����F'r�CB��D��]�!���!�!k٭b&o�hϿ]̬%�������9�(U���h���8�q�6�{5�&�2�jXV�`��������O)P�8��?��R�D��>M�k��[��A�s@�[�*��:>]p:�C�3Ul$@xK�;+�Wnh��0��~�.���y�0�+hE&C܍�Y#�i!%TJ���c�UADb�~H��N	����������@ �R䆍 [�SW)^�*A%V�*�gh\f�&�VG���Mqs�k��Z��E��7ũؤ�Vqs`g]C���	���t���o�.ڿv%�""&6��Q�o���|~�E!"�XR4
ϋ�X
R�9�s�:�kk���h�5���s>b��X�� |O$�b��(�E��$ϥ.:&I�
}y�(nB��ک��5��x{]7LXNcM�z\�<$f�	h��jT��)'���R�"9��mA&(��0?|�;��w��-�%�/O`���z1�J/�k���N��sn%r�N��& F����7����Fr��8%��������5�v,=�Ṭ;�},'&`�|��Te!�o�Z���5�[�� �A�ە]�憡J\��	�N�+ZDj����R9����O�,'@�{�Q��:q͌���8vd�.[�a����4�i��9b�q�i�?E�7^ʎ�O	�M�|ܨ.�>k�����-��J�Mޟ2�A��e�W��n���i���@�Ĵ���
ձ�S��]"�x��W	w`��-��n=Bn�Gnf;�db�ƹ�?��¾�־S%^�@ ��;�W�ɇ��)�N����%���x��}��p�C�	�~i̶�BK�����R�l�����	�Q���Z���_�+E4��'�^B�j�d�PK�^Z���Q=�1\8Eؤ.&��1!���{c��z*���r����{��7yȰ���^���%��'�����|����m�3��@���J��mbQ鉅�:fG��$��#\EF������u�ۧ�4�~,��5R*�ӊs;x�촮�ݺ�����ޘ}�۲A�Ly�N�&�fd�g1С")#2=n[è�̇1?��La��?��A�z���5�������d�Yg���[�]9\�����������=A�~���I�G~s��42����g־������Sٰ2�~�)_R����F�`��wn�1+��8��KT~{bc��G|�4+�xE=��z�C}��j���X� ��2������ĉ04�~��Wږ�/VW*���45��5�+���A5�������J����r�D�ju�'N�[N����Y	)��_�՚�׿p�����AQs��V)t��]�)�F �����m��@�A��;I�1���HK9��1I?َL��!���t\h)t�WH�f.�4?}i$LY�8N�U5���3C������1⢝Ճ�oK���MC�O���5��Q�m��8�fZh�@P��P�Y��=C������C77u��౽�d:���v�k�!3�O�|����n�*Z2�����|&�Tjq7��)��߯��6&.�5���_:�?�C^Q�`aI��T�ˍ�{��ڞ���q4H5��L�87gP,�����P�9��@R�ѥ�@*��������n�Ξ\�y�;��%��u����"������_�2Y�w@ 9V�6��A�[��y�%�DF�]�:�4��ç!�:���Y1��S{��4��g�OY��w����TD�:��Bz�C�;ox`�Vq漉X�V@��Ƹ��qo]��P(G`aۘ���B��&�Ȇ����5O*���2P$�Q>ɗW�r���C�Q�)�A���^���6���۹{C�'�T�t���d<�pGe�* ��>�l��F7�}�<����L٭��Ѻ��j�4]�����Q�����?��
O���[v�)�7���%&�1&��)�2�:�L�F �H�F�\<_B��k ~����o�B����F��(���W�//-�Z��㾘Am�L��������F��iܗ�Z����	�&N�U[�AV�*�����b�D` p]h����j ?2��S|�^������'a�:�9��wV��=/��,;¦����%�������OoG��K^�u�F�ʶ��G�G/����;�/�̀;	��w�S����Yo�k+�-�}�k�s�a��m��t�����˕���@�k��3m��qтr���R�B�$��(٥��
P���]B�N �nm���n�qL�4�VI�!��S���mn&�]\x�9��6�`�A�qT�#%��֥�U*S2[�%X����=X�HF�� ��z-2������=������ހ��Uߋ�^�9��DwD[|=3�@��~�D�U��"x��Yc������xJ�-lV�!\�]g(Ld�\n#aN�Sl���*��*�)�~�;��?�tI?'iK8���#�Ub<\u��f�
 D�^��i�'`��+KV���S�������"H5�y��B�1gƘ�JI��֎5�	���!����|���Q��tn�!4
���e"(����<�)���"�T�_���_ik�[�M��7UI����Ɣ5�Ny �Pw�V)�[i�%$o�t�Xl	°n���)@�s�\��">YBY�	���o.��R��R y����ivV�o�p5?�tqj��R��w$�QP�ƸJ�:����D�����L����8ېu
�iLV	��cpe��u$�� ������=.w?�L�qu������L`�<�݇����F|��u�ח���iL���?�ٹx�m6S�Ι��f����U8<�c���p/rMׅ�r��������탇Jon��
�_�K��i�t�"�������=Y.�N劉�+1(��XH@�j�<\ǹW֏��w|~
?s���L���_���LGN�bZd/���Kuִ�S� ��/��싶q���Znj��]�<����p��$?>`8��������6���I�f�37�����hmRYF�Yߪ��RZW�a�x�Fd�{-��Z�_S���� ��g��$O�CY�*�:AiHz��F��s���̈́�t,y/-߳l_��L����_�vw��>QJ�$�D������A��X׃��W��5��Α9��W��jA��j���ӗ+�Y�J �(�v���\r����$o���=dL��:4r�#��$ٽ�o��9�O^�5�q�w-ߋ��{;�w'�Bpץ��}��h�>k�:]��:�dn2s�P*!�E�=�����X����=ߝ9<5�3�0��������{��r�ޫ�ћǯ).�c���ɋ4��hhG��N�Dr*��������"������0.��ߓ���n&��k*�C�E��w�	�A{�;�4ڙ;��ZLNYu��떵'߫����R���<m�,���r�Km�M�[�'�З�F^�+vY��4�����$�"�uDJ�J�҅~�B���z�}�xY���<����r��e�%b���KɢB���(�>;xݵ��UT��>xNd��Ҵ�iJXE��T���>{bCn��?\X�^����i�]����\�X[�-pr2�B������*�f*�}�v�w
�/�����AL�oџ����i=����88��T_��A��j�i+�@bO����X7��m/��F<j�MJGMY�sz]dg�l������$`�A�S����d��`$TŒ|#�+�t�x���P9	�u�'�ӟ�UT�1�C؋�qhĤV~,PH>(w���&�dKИd��%�o��~�K5���$4���|�t�����*T]���������56A�(1��Bi�`d���U��×�9�Fgm�e㱴G�����u�Ssh3��O�_U����X�v�j����]������o�<�;h|��	����*Ni�e�O`	/� �ǜ����gO|�E|��y0�)l'�\�
8�O�&=�)��l�h}�k���f��E%�z&4���Zĳ�Ӵ�6=`�ޡ0���B��{�3�yXJ�>�e�s��|{1��Ǩ�?@���r��/�⻎1�O�(�GW7�;f��[e�H�~)o���r>�N8�x]�}2�!��~�S��c_E{P*��3�'�ڐ��ox�M#컑���m�W�=�1���Q0�ZȘ1h�o|u�xhyV*��6ޝ�t�l�(�����Q(@[<S���sl���&�d苏G��"���2�� ��<x rh� �����ꥊ����<�RV�:�@G��u С�3 �	��.h��j4䉬�k�0�_�t�u����4���]��zX[T����G}XC @
4s3�+��V)��~$���d����>L�:�)(��R%����E����K�U\D���S�����8��P����cg��`h Ih���'a����5��ȿ�I�:�ey*�� R/DŨ�7�
������"6'E;�j��]�p�4	mw�e�E]W��(��^���Ԑxr�[ D�x�7���{ȋ:zA�rJ2�v޳�|�w�����u4B��K�dN��E1)p�s&�O8ϡ��	siL��V�v�>穥�s}\��F�|cjSr���W~��G�p��-*t)N�f��Uo�ϋ.����g�uRN�PT��M��F�����,�5O�/�i'��6c|��Y��(D�r&��,�R ��;�3��*7�0�D+h�0�h�`��0:O�.�
R�	F���sp|��R#]�@N��r>�U��*�8���y�gXC
Y���V�} ��tK$�����e��F(S��߭^�����F��c��Xi΍N�Q�"8�/�{��� �d�����(��;�/b5��8�y�TC.+B�f����Z�MK�O�T2ʤ�b�ѐ�Ü��0o�m�rG������~���:�;��.�F��w!����,���H.�&}��Y�:�o9�V�\Ӏa�f��[9�m)t�o��]σ��@����CD���wYXRK^�7��qe����2���xyv��Qe�qY�ڭV�K?Ga�o����������CÚ���p�	�<��0��/��B0O�A�BT;r�����jR ղoT���j��.�!��l�E��l16#��>z�%{�4��ۃ��_A�����lm���;�^h�OY~vǉ:��p��,Lp�
`��7?�B�NA&*}寮��R��)QJ���G����x���{�v���ر�Nd��4.���v�m��"�^ɷDrV�c���i�D��3�獻�G���@dY��)��Ƚ(;�C�s�2zo3��wt�z'�8��0X%j�ٞ�f�
e��D�
�|P�$���8,���)E7����Κ������r::���s�c�\�de/�,����a�Ċ�[xt��o���}qda¤����C����%�_ĩ��5�q]�0�R�vS�-����[N�E��L�y�~I���5��K��N���W�����e�)�'�a(%]INQ�5NVs�\㗳�W;��^��i�J\aɰ�(�0��̋��[���:�/�T�)�
'�T}��K�{7H�;�����]0	��B��к���*�Gtq�-�c0���%S�/�^Ѫm��!�*K[��U�CU��3�g���SW:)ilV�5���r,DC�|t�(;��"�JyF�q�TD�EP�9�ۘ�@U����V�3-V���'���^�tpԴ.6;� ���`iB\��g�o)4pOm�<�3)�<�k>$��EK����"#�;k[�)���۾�BnX9x@̽����r��J�4q��uv�?��mq%���؝�8�ry����I�9� c<ө� �xQ�0���oِ�����P4�]�v�$�;8�i�DIGU����3�,��E*��ҡ��>;�����K���y��*6J �b�pJ)�.	
�g˳��9j��}�:�1�(K��W2�Ɩ@YPsL�]��B���d�4����7����`�A<�zH�J�=�p���(�i�DÜe�!��7�&�g������a�ç5@Z)��A�U=�C��>Ճ�֣닅!d]16���Ɏ8ja�<��A� ���bCX�:.��ô�<�6�a�0���o�/2�^X\��W3DN���a(��$�͕0��P	%ݴ��݋S����M�SA�;d�z�Z�������{��ߧ�bT���UO�+��[�L*�v=5��g6�e�@9��Zk3�m������!�x�GW6$V�	�4=��a�5GxE����P��۰�fkZ�T]�y�3��@����� ���f�s��oR�t���9�wLP�cwcG��!Ti�4�����^�/�d���Ф��A̚�F�.���=�<����o��˽d��dg�CC��}�G�P�p���{� Z������9�X���&��+Z��+1?�\�V�����HBsn^~�qz<c�)����n���|�[ �t���(H�f�U"^V�A��cu���|\jv��<z\li&�$�ґ��|8/7e���"�w���k}˘�R��*���h�7�jlu��a�Ѹ�JiN���S	���Н5C? Ǿ�� ,�I(��y���p�P�f�ˎ���s�����	��BI)'�o����A�xihz���M�8}�U_5d[�vO���f�x��1q�u92���Z?��
��81���ސ�����W�N��)��n7W��B�F������!��$\uڱ���z�S��kڿ+�ݓ?yOOC�q��ΤG���Ĉ�c��R�w�H{�f�$���#V.~� :���C,P?�{]G�<�^	��Bo��0E�"��2�#��N5��l���x�-��}��T�'��W��&Y5��j�Z��5XӴ��f�bu7p�.�,��hZkE��6�n=��i4������!�)|A,Y�s����P�O�Ry��1�n$2�{C�Jm�*�5��o-��={��1��ӽ:Լ$�S�D
HV�fYs�Y�U�w�y;������2qQ�ȴO
�Y��H.@F?֓>ο,p��H�/-w؎	��鞣#?�k<1 �,�w�en{.s�,T�%� '��J�&��'GN\�mX�t
�14\اmYl�y�:��b�5	�Rg0�7�6 �9��	�Y��h�F�-���}�
��O�K�lZP	'3���.�`Tu�Ͷ)NՏL
c�ct>t�����x|��*B��V�k�W-S#Bc�h.��i������P��e�\$�ꌐ/1&�?��y���2�t�k�IۭEWȌw(<g`��P�aq�l�m'g�<~���*��A.�7�|�-�� �m[��Ng�rt�;���	�h�t���=}�l��P.1� ���
ZMH�-jx��T�i`U#�"~���?�Ș��8���E+�ގ�(����eVq�r�7S?�|&�Sd;딘�z)k�P=ӛ �j��"��������?~v�����Xag=,cs�ż��C�ɝ�+�q�qb�NB�k�N��#<��`�A��<��q?�,������`��Zt�[��ؘ�>���C �����L��*sUU-�tp�%k�<|�_>���!����B��֏�_|ǻhx_�U݆���d�ڧiT�V�)^d�w��"'�r� ���LQ��[�5��Z�ΑJ�x��_=c�<4G���T�a��ȼ����tI-�S��M?"�q�
(e�c:ewʴ1��.yg�0_��R-b�wZ*��[��>�\"����G>�M��n��.��X��)��0[�?ka��H�b��i���kdx���,�R}��ߓ�)�xq]�x�0��}W��)�����Dg��*��̺_`~S�T�_�Q]+���R@�7�9�ދ���{�����RGQ��[��eI��#�
(�����Bjl�,�,�e�ɕ����Д����� �¬v<�4�T��uYc�^��B�����q��a��8d��.�:;�a��◓�5�1�jO"�!��O��K����A�`=�����@~�
����Y���=>\ҭ@ŕ�K�sԇ�sn�^p���y8{��T���b
M&klwY.��q�p���"3����c6o̚�����i�K����U;E���-��"��3{�a�������ʟ_��ؤl�񼛈����VTs>8�w�2�Z��I 'l2���@��F:��E���d%ӏ�;s;U��x>.XƮ�.��,�{^�H��j��X1�#c1J��+�ɹ��KAPA�M��S�~����U'���,1� ��{�e������N}ҽˑ�#����m�r'|��]m�$���g��t��Yh8A�[O%���P܅	&Ǽ��V|�"O!K�K_��0,�NH�{Q�/U?ɓ���TeɌ({���H��"�C|�gm���J��m���ch��4�q�e$�>�D�N��9㻖I$|�h��ċX<�L�$;�ny�*�f$�6���A.?�@*՝�sC�ڴX���L�PQm�������is��x��yWM?SF.oD�*��� P#�xo\I��*��J���'�@D�^O��f׿+����ԍ�E㗌��j�'��H,����YVl�n� \p2s���*H���P�y7p:�?��M������-<u�:��أ�J8%����a��>�<�Ӽ{	,OH�#�'�$2F/��;���Hwq����w-�G:&�A\�_ۿ�Đ��YE���[�,��+4�A�S#K��U8�NE[����n�\1�/Y��?f)�s�$����+���ٞ�r�e ��ڹ�9��������{3��G6(��	nH��L�:��A؀I@�A&'�^qݶ���=��k���r���;4Q ��
�q^�\���b7��v�%�\M�u��+���h��vB�W��).����?V_�-]�@�.�(���U٭���.>����	N[j�I�y���ф��o{���Y��>������Yq��"I{�� �b'��Ǹs	2�|��G�+KK4PZa��3Hu�fg�ו�!Va5K��a�S���ҰM�#��'|�+�P�l)����Zޙl��m ������G��7�����A�5��H<s�0�����H���?��;����e�"������_��e����!臒���K��sF�f�W�Ƶ$�S�>��(^�L=��{?RYZ>�F���> ��O�?�2$̀�I�z��t�x�Gt�İ��ׄݓ"�4S������6��lQĨ1�o��Ir��ra�����7����������Ed��+�b]vJep���дSc+]P0h��G�R�?%� h"S3�G���E�Z�V�hRވ�EZ�*D�[���Em3F]��/PF{�;6��W@�Çq�7.�e:Lw?7K���-�ކO����|K̅zg�<���@��%⽝��В�Gf�w�N*'���I�DHb��"V��6j>KC_J�H�	�������ǝ2�e�m����� i_�,²np
�덢l48h���H���(FݣM�S��}e�cT���hwF6�<���A'
�ڤ��u�Jg,��L'-���k��Jm�!�N��������m�.��D�?ܳb�L�\��vB�r�R�y|K��*���$?�[de��ؔ�aS�~ �F�aZ�md;���(|R�M%C���뉩�J�.����7�75�Y���ܞ���C����t�ѱPԸ���;{������jZV���DٖF������9V�e6���V��q�K �rN���u��ޅ7�E1��C��#����_�s�7_�`AQ�v(5%�S�P��K�}7� H�O����q����1�t7��e tF��f�]�Dy�{�RJ-�U��z�3���������((��l���n���4��%)�Β�6�OܳG��d	�JKO��+���S��_"Vp�B��7ܴ�Y�Fp^	k\�{������ �ps�♌�Zws��%:TD�2���h۠*3��?>����E�S�-��8�z�b-�WR�>3Q�%���c�I������lVĊ�]��OK��\��&6��;�v���{YoL��"�o���p���ąǠ�ްh�m��o|{[�i@8�������?�g�q����i;��x���~�u�b�;�-E�"b**�pl_����I}6�x�)Á�U�DY��狶�c��3�Z
��z�/p43��83 �����2���_d�Xƴ8���LQf��|֛�8�8Ss���u�s���pP�'��# ȉۜM�ny;�����
�G�ճ����mU�}���C)b���P!��ڰr_Au���NI��<9��Z��0�ޖq�Vm�r�dţ��>�T:4�>6[�:�q����,��0e��YE&�������Q���V��ߙ˨�Ƴ��ù���G4J?p� �	��Y��� f�ΉYkvTW�4���K��9ÊI��y΍�?΀3��x�d@T`T!�)�X[�,�.����|�㱜��<LW�	�jGP�ٜC��y��Y�m��G��=(�o���t(����:�V��2���zr3��j��O2@m��O��������i�=�
}�J��Ar�hHx�dz�g�WGeA�JQ�����<zbҧ9�Lvr]wi��l�˪sw�x@�?�������.MS�,���b׹$/Ë�QW��o�y6���Â����xe��)s���m���o��y>�ʵ�#).�W�8_��)�D*�]�\��M.�ծ��m�3�O�8[U�3�!G׭�H��w,�>�b��D*�,�{�HT���)2.NS+�RT�	3#�����QM��h!�G{o��_8�f(ۤP��=Oubi�&�tY�KB�s�F��cJi�&��6���6+�[?�\^k�c/r;d]��Y5�W��������ͨ@���~�� �&�!BI���M���'ȿFiڑ�2�ζ�0�S��g&Zї_�"���;aj&/áIBq��Wg(+�gٟ㮓��ڡB���i}�!5N28'�n{�am�9�9w��]Wqx�����j�I�O��䕵�mZl�����'�.d�
ۙ��+���9��/@`����A��r�Y��ĳH|�	LЗ��p�L��ak�w����@�0�!���ᮕ��/��z�*��������>��
�<c~:pq�A�JA�G&�w�@.���dzI��ޞe�c^#��v��M��ϧ�Xn(t+\H���[_?9J��F(�'�;���'��9]�g��Z�Q��[�L�M��8W]�o+�vm�i'��e��v��F]q3���&{K�� j;m�l��$��OΗ&�vz�+4U�WT`̯r��crKsE?u
����v�1g��J1
ml:�g1̚�\�Rv�;��X��0���т���U�zʁ{��8	p(���.��9�Cs��{Ք�I2����U��uµw�T�A扣�>0�w�s�	}E���᫭�X�����(���֒O�5�2�	��W���l{�I2h�D��+q��RM�:ԉ'�n�`�B#�n�T	;�Sj-�/Iޕ�d�(�/�f��"���m���3��ĵ�����T,�H#Ş�����bDi�?�%W>��lA7�����j������z�h�r��nK֎��!e 8%I�]��^M�<��EV��(�F���I������vƵU!�Ԋd<�ck���V�w�*���r>Eꡅ�@�
�DB'E���P��0{jh%�f@�Ev�e�=��i��7�D�r����ەڂ�vYGRQ�����dfL�/�	������ѬV3�t��-��E�Vfy�`C��� *�c���rq����%���! �+tS����9� U�d��xX=I1}�*f�D��Ӈ+�zi��A�R�(ڑdfs�_��E�]��,YyrJd'��rͻ��$9zOq��^��9	�e�D�I�L�fl|yF�UT�I���E��f��.���$\�>��p#�w�]�
������B�ws�4����xT�y W��f�Ƀib���1β#X��� �V7�&4�HC7XL�b�F�k�9y;��>%bv��$*c�f��&=�=%�[�8�>X���fɸ�y�~ʂh�]��S�S6�\�п	#�&0�u��bmº9�?C�5<�1����]̭�AD�y}m_�9`����Hl�QA�9,��W%�e��J~xH5��@�΋�����vaj��A���b��R�Ӗơ�؉#�H'�ɻ�`I��	OjMI��˕9�Q=���O�6�.Z�yNg���GY2���I�1������r���*�HC��GK�[T� x�Ү���	�x��)�����q���S����N��_<�ه!���r�F���:���
�ň�1ĂOŦ�M���i�0�rD�w4�
�F�&n���*W��x8k��Y��n�v�.�Xս���B��86�=�*�;�i���
�<>X��@SI�����u,���F��j�}� �^[	�����i'����d�+Y\{߫�M����D�b�gk��0�͵/U��	��� �%���k����9^7�Wj�镭 �X>tnV�(��v��w!v�N[�'ӟ:pa��EUݾ������߱�w�I��h��o�u8z}�>���o@��˨�,�8�^Y��u�l����Z�#���zP?�X��4��M5SU��M�F���y��p�T�7��~s/�r���T���$Wdtt3�L��Q�:={A�� t���g
��+2���	��8�4�������!?M�6b�du?ZC��Ų��x� �LZ�	}�
�bA�A+q��B�M�QBc�D��`!�G-	��?�\gQ�� "�����F3d�r��(��CW�D���p����!L (
֩���*B*��d�(�_�Q��h�A�xL�\|���_��f3ߘ5�c�򎄫G-��h�VU@c���l?�bx+�X�ר쬐���ʚTރ-0��[��NÔ��h�iTBX�ވ�b�戇Pz=��V��u:�)�X�o�ދ������Xl=��h�]�4g|g+�dY���.�Bqy�+Ր�������ھ�R���F�.���
B&�6���z��)6@ޏ�#o�� �88�eEŽ��݉�[~xuPo}��E���,B�C�� V(�^?���*-W]�N�/H`��w���ڈ�vGp~!'7�e� ��m���5�<���8%�B��4C�{~ݯ,$��6{~0�Q͛�'��k���֚%�0�K�j�!,�7	�'!�j#��9�{"�z[&��F2���j�"q+�]�{B�j�K����-�#M����������i��Hf6i�d����	��)Ĳ��Y�����o�����,��9;�p��Pu������3�&P���o�B�����=s~���Sr�Y��<
�4�U1_�%a=P�I�� ��o�e�a(�ӝ��A�C���=�����Q�c����fr|�0�����'E�|N0��W���=֠Y���YV���^�X��v�7�B�9)@R$��Ė�e�bM���t8i/)l|�g�"s���SH�F�eU�����3�ee��K��7�]��w���C�MD$`ү1���,�ߪ�K!� u��~g�8��]�	"�w���*��
4��X{(�).TX�X��h�Pg�)�϶�����]��yn�@;2�Z�9��"��ķ8o2�=<l-�C�-ǉ�����!z�WOl��I�I��Ӧ�x�o����(d��#y��wO�����1�I#���	<�d��D��{��`��S�6�2�h����j�!N)AD��ðA>\����Ĕ�FW`���6�
���T�`�
��Z��=�^�T����L����R"����#��1C'�r��CYBPV�hW�s��z/�3��z>O�g�@���3T�����1�
۷u���ܦ�$g8-��:Շp���!."Uch��A���׾�q��6S�A�q���F����g��-:��19A����y�����E���1'wפ��ǹ�)s�wN�u.+I6=&�lQ̒�0O7S��h⟘@>�CtȖ��Ӽ�v�s�r+���[��~�������Bo���k�6�j�d�=zEA��YQ-�B�^�b1j��߲k#~��|���Y{Г(�Q��Թ�F�x�L��٘L3�fmݙ!S�?'��9:ovk��!�)�Gw_������׉�����Þ͍��U�OMFt�sF�x)٭ѷ\����0��k�n%��6����[2�=<��6I,�<��N��t����>�מ`�;7�u^u:�\�i)�p�Ͽ��}������,8_�a]ۋ1K�7� ����ښAS���g�>9z-�3)hE�L�0���K_�&���̜�[Ï�uc�(��M�CU_C.=h��Nzв�'}�O8�u^j�q�P���ܽ�s���ba{$u���K��R�G����~��S����/_���x2ʳBb�+*������ky�Q?T��Pq|��S������� 9ֶ��K/BY�, Q�}������E��O�'�M��F;	\Z��x1�P
���g5��u�&�&�[�+�qޠ�
n��-ꐐH����1<<A�_��qB������҄.�y3m�'�î��m���;_]ːlm�)��.��������E�u:�s$����<��72�GQT"w���n�dy�����D�a��A��iV�%�h6�|1����3a ���/�}�w����V��Aq��$�z(�-�iK�/nó��N�@U���8~��xR���\I�vO*�.�������,�"��;���6�+h���4�m���s���=��fI7�e�r�u�Yԩأ-H'������N�[x�GF�oM�튶�g[>��i�J˙̷gM�zj#��Ws���r�4�JTwTc������i�����,��0J�D���2�3�9Z3�>��qYi��h9V�3B-w��&�-�=qV;�V�������P�(��KO��׋TH��H�fa��:t�b~gZ��E\�0�N��J�6n)��|5Ql�/gqT2IC�sHt�l,�� ���N0�L�	5$K^��l�!ű)���d��}�EPe$�4�ה^!\�Y7���d���/��*��8p�֊�һ�(���Ҿw5J(Ď�y�|SeAUH%��@��"�����m��\����R��|��%�= VCkV����q��4�qܞ��!C��	�(�K������f�Y�G���UĽ�wy��@,\��A�Tʖ�S?�~��Ҍ���6�C(N}��t��vRp)����.OG�6ַ�^�b�1�����ɂ�C^,�0i�hesV0�R�Ң��ʾf�j�pqyayZ�6g��̪�^(f��/}��8�ov�8��`�h��@&a9�T"���ֵ�w@��;̦��Qi.�yYY�D~�ʕ�96=!I�l{�,>1��#vCv�IYԹ9�c\.o�ȁ�y����е���U�Q����-���}a�$7��Fs5��U:�i��~�y��@d�*D�AP.�(�G%f@�As6�w<)�F?�1�c��G&.���50t ���䚼1J08:ױz=���S�9H[�`E>�rN��p1�N���%2�{���J�����'�>L�/�aR��|n;U�92��k?��b��Z�>�^���Lz4_��|��V��$	������y�7���ܕ��R��M�՘*�Uk�t�>�a�M�}�OQ��}H}~t~��`<Z�cQ/�z�Pq���}�G,ٟ��#���O5�ܬRa��}���8n����՞6i6�1�S���߁��!,A7I���8p��9�/���|ۗ�mi�?|� ~U��94�h{�^�z1�)������k���jzy�#H�H�/q�t��E��Y�rwP�S-pk1��D{���嵥�?<"�n�x^���@��f���儒8���QPeZES-�1~� tPe�؆��%-�h꣼�7H�g�(�ܟ�S���N�E��轵��{��,uVtx�ojcV���H�<m�kMR��F�+�B�m��;]53%�5�tsE��\�U�}Aݣ)�1ףlM��Cmf�悪 ^!�.K�rN;�R��۽�%�gD�2����PH-/��5'�b��f����0E���c�q��.��YL(f�h�2���gU��T�F�P�����/�8?�i�@�Ν�OlYH`7���|ˣ���!GbOyH��6<l��[��r�|�שˋ�C_�>��ǎg������]�/*��N<�ޒ%1��q-��,El���Dӳ�*d����/^8���	�ׁ�)o�-"�o�(���,^��լ�B�Ա�>H�r8O�-�J����=Y��=%��wW@_�.!�Z�����nk�J8�;I�6��"�}ǎn'3�$� ��&̀�P�'S{d�n���$��	�j��QE��5���|�l��(�! w���H୵���YIЩ��ۇP�&�̿`�ެX�}|�$��O����ܿ^�y��h��#����t�a91���(K-�w=����^���ѐ/��*vZ�kv�Ԗ��̫�̅w��ރ4��Џ$��kH��7��犃 �.�(ZÓF�l`y���60�6��chr��5��#�p�x �<�$V���Y��pEK��`S����ٚ1����Q"���I���]Ӎ�ͫ�y�����XTo�K5k�3�y�{HpDɞ��,���l��@E`
|A�H��7)h^{�Y܎�.�W��.��]���!.1�����+6���)�P�Y2ML܄��=��,�����$�и�B�z��]Sǈ,K	��?L`�X���z�Z`�ҵ��{����.���Uu�"q}��"~��ײ�B�� �eM��|�g��9�l:h�Me���w�T����L�s'ǹ�p�$"�fӰ��jc���#8>a}x?��5�7�<v'�)��&��}A�� *V�8����.�]�n�'����~:`L�D����V`2B�bÑ�}�Ws9'�fr��&zJ�q�Fؖ��"��O�����e�uհMNM%9&֞������m֥�;�����'���.�.-G�S,��C��+��r_��]��/!�\��3:xАbg���Z.�F�#���e֑���Y,�7�Da0���^�)j 595�ļ��o�s���qV����-�l�>��a�X��|�k��W�S������I��E�)��wA��>��Z� �E���[6�r*V����<�K�%�Fm$��ZM�t�iݷj�wv�T�������h���۩��e��g[:h|@6㲯���&��SSC�u���J��Ly`�coFn� bYJ���-��w�l�
��/kYW#FA���v�"�=��M)�o �~��Ύvk0sv��dM֔<;�u-CS�Eª��%�K\}�~m\D��e�� ����2?ݑ������!ʿ-���ZA�T#��@&�06��N'�������v���i4Q�� 2,\����5�����1�-.쥞ݼg�^&U^R�f�G|z}��/hp�f��9�h�t�mK9�db��=\�W��$�����E�9
K�w�W�����7����I�CG�m=H��h%��tS5�b�/��h�u#�/���Т����W��t�������`M�y����7ڞQ(� [_���\\smP���ӻ�3�:�U����.��*�����+���%{H�������CDpz{U�	?��-W�EP�z9��q��<� �Sp�*�u+�+���ܮ��4��3��L3�.�>)%�k+�w�14>}�ެ4��K3���Ki���;�6+�	g�I�[�1��a�.��~BKe�CW�� ;�O3������=���0���v^��\u��}�������	,C	���@�Ԏ�e��4��Q��b�����r�z�5|P�FƆ'����^����������)��"�)�P9�����t���~a�mC]�`�+�P�g����,���*�M+?�h2졗i��̍� G��J�1;fS�O�$����(х��j��i-A��KTc�B��O�v`@,�D#��:���/�Я�$�t��^���'�H$
s��^HVu|1�@e�&�d���Y$�{��v�]m��#��O�:6���hV�d��m���<�0Q����3uUv�m���.齇�Rx�����,�wG(��h�g�ʡ�R�j��/���vM��6��ޘ7ys֑�����k%�,e%�b�;��T/��[9��|Ƴ!�]�fTuN#h 9]��n%�"h�=�h�oZl$`�s����q@\�Y �qI�Nn�P,�!yv�����_�t2��x�}�U|zbq�ut���[���n\��F��P����{��k�
BN�#��8�.��vG�r�_-���!�La�$=U>$�)�0�?G���3B@�ޔՕk~lF���z��n�%mQ�@Hrk��-��YӚ$.�8�F�jW����W(z-�[��O�y��Y}(X��}o[��]1��`�X�����_��@�}z��=�Fg��e虦�$�;�o�DP���{πXq,a�WO�c�eQ-4�I���\U�����<	iKݡ�Z��,�[OJ�Z����/�;\�>S�~����rLMّ3�_�����sD*BF�b��J34�N�=Ep�����F��u[x���y8lw���-|4V�CQ�G%I�a#D����E=�tl�U$�cu���;���>#�v@	�p�X�'�5��>M~7���!mP�P��z7��ưΊ��`���dY���#�H�1d��S�Gg�B_�3��M Xa(���Wj���tI��nQ�����w��WЌ����kne��|")O��<9��J���/��!x��5��FfkY�"d���g�5��uGE<Z29ff�g|���5}�_�X�J9?<!��ȥ|�NE��?ׄuiuD!�LTZ �D�;v��	�B����92ݶF��-���+�����^��J0���-�g��ȭ�7̪Z"��xBzs>M�%��"	s������c��A�E)�(�
�_���4;��'#����K"h�9��+�l�`zm����@�+�1ϴ�oDe��/�w<-�'�A	��q��*���|�&X�)��w�:��@h�V3բ
A�0.��ʥ���5�x�-�n��tnv�w�=:L�q:��95)��@��A�K�V��$��Md��Y��=����xT�U�)��Q#�"h��CLCpxnHH�N{N�9��/ Pk�i�i˲�=�x�R �X��4p#��*�ܿE���r����K��]����t�~:1�k�Z�$p��������F�ʎ��gž>!��3Q�l�����7� HsF�낰�[n�WgJ%��m��J�A����Q���_��9�U��Qk�Nɻ�F�,�'�0�m'���!�ʹ��� =9~r��P�P?�n�2��&nY������16�z�m"������?�?����m�F�+��	�B�J�R��,�᥎e�d@�1����z����%�	���
�����e���L���-$�f��~���A�Y��5	���K�M��)��c��F��s�^�U�wɷ���|fD�},+߳�$��^�Z�&m9�ߩ&mL�&A��;S�پ�dߧ�!{3?�G2]�C���5��?�qn�`G��q'E�СTՃ��*��	+y�J�El�_�� ޶g����)(�e��h�>4�� Y���.8�)�4$��?�����Ĩ�
�>�o�>��:+�g�͕D;(��bjl+ Ȩ̋�7�P�Ur���_������T.Aт�`c���8�Y\�H���̌�ґ7��_�,̢��h�P��z.��k!(p1܈-L�F����zKó��Ӣ���z}G�.�vP��,߮n:�5B�G�;�n	������t1��.xB-���V�޶܃{٪X��ֶ@,�T�s����2F/��f�bK#�)�^�fF8�Z�t��^�46~j�����@զ$�$Hni���\�t[�;ؖ���W}YH�����5�cAf�9��䕫���P��T(�v���}bB���B��BV��MFG:����٠pɥ���7J�������Rު�YNq�E�uy�nw4x�۹�`���4� �Q����KN'I�o�DXz�Sc�e��u�"��ҝF�n�'n�/����� ?V]	b�oX�-�Ej��l���j_���ܕ�G���ݵ���)s�N|h]f)T~�KQ�ؐ+Ŗ�o�L���.J_2��������;��#��B�F!�Ƣ���!����Sߑ47 AT��.�i�����u���dN��X�[#��u��7uɟ��xBŽ4�	�_���!��'�}�R`�L�w�)l��V���b��K�����ѣ�.��崦�)����o�M�0�F5q�1HU��,4��^�b?�y�������i��P��oƧ��m:=��mG5�?*��l�I�'<��
_�I���}2v8p <��`h2����x#� IO��FF��dc�SO���us�������T�{�U2�ɽ��b�ҡ^��YO~�����1���4j:~RQ×J�U"��R�cN��QXB�[*�����e��&4Q�YCj��tT}R��"�4�����5$C;ZgJ�I���؄Nd�qg��l����"�����,����R:L��el��6��R=���S+�>��1�>Pm�<��KT��"d�ᴌ7����{� �V��R	:M9v�Mػ���A��^����Σ| ��Eb�6X�%%倝Qw=(�x�9�X/���o�&�*�"���{�	�l�-Σ&v�B�Tp���lR;vI�[�OV�N�����v��P�C/Y�~�w�Kꊓ��r64lD�QqH����"��nSok r��a����0HVM��,8332{pр\L��3�I�xD1u�lU�z���;��íEU�"��IV���"�׍/�n^��B*<�Q�:v�	�Z<ׇ����g������(��-�`�E��P��{���jD�
��f�fh�����{�+����t�y�2BWq��p
���c�s��8Q�~����ֹa�Lc2���Hޥ�kﶏQ��Sd�R�Bni�Vi����ӑs��]dZv��ݲ'��fx^h�N�:�
������^��ɹ�ٞ,�a��=;y�X�zt,�S!W𥔓��QR�&�w����2�v'EU���H�a����.i1����rOR�Tӛ���MҠV6	&���ʧ��I.�TcZ����Y�~�SR�'[�:+�e�0��T�yפ4�#�yI=?�r��,̧�E���QykVa$G4�ڦ���Ҡ�6��M�1L�=��i(���K�}N����<L��"JNg,��q�qΡ�������#%l��0��Կg�\�4]L!��&� �'+�����1_���9��N�$�*�F�|}:�=����kj��ܮCG��b�˪���V�A��-B�'u��e �\?=R7�d�/��c&|'���h�-I��?�g�GF���⯨3
�� ��'��:]ޡ�[/͊	��I�}!P��x!�$k��!ý9����E��JB#@FĪ���Q�7ܿM�q����;�s�q���]�H�O�V"?Bq�-�����&	o��L��o(���9e��o�*�u�w}SR�-uC��FT���H�f�X��ka�2�g��=�N=����zT�+y��e1枋[�d����=���5d�U5��-K���m8�+��Bqɜ"o�l�䦨̱�>���Eg(C�������t�#�J��j�L��du�� ��շPF�C�4��PyL+<	 �I��}�#��=b����T1�vms����n2�[�Zn%���w(��f�(��ȫB�7�j�Ƥ�O��f8�����|޵x��6���-��k�[�:�@9)r�!����4ՙ�'���'����p�1���hPIglR����.�ϔ���䏢J��@L�i��RXE�������}�tF�½͂�8u~�E�6Lw׻ �'*|a������h#�ܗ�.����/���#���;Hz�#H" ��Ʉ	>`u�H���5�>�=\K;M3E�c�����j��s7<[����6N��Ț	y�$
s�o���L�����p�ӎ�Έ.{��]�"��
eTzMH`/�셹�2O@�U��Pu��<
�Ƞ��T����ٞ����B(�����2��a+|>�#=��c׃��\���j�<)�ᨚ�RwVs�kT����"�W8� Ȟ�L~$���iZB��=���A.����
��q����Yfw佱�Ɯ���uC�q�S?T 6Ni�	��'�{�,ï[Kd(����=q_����_�>c�&X�QT���]�q�N��g��Su�]��w��{������4��4�M�z��!��[�ڮK,�o�e�Ee��I�v?@y!̰i*,ah�M4n�.cz�:F;�%H!�o`�@���AԗBۈ�_��� M$\Jm�gl:]%�Yt-����MOs�k~��F�T�Z�%[��y���_�v��E��O��b��<ɢm��2�?R6׿Y&�:4"�`.&��t��sbK��?�7R����ҝ�+4��T:,�i��/MY������f]>�7��ȂI�J��-2'e:�%Hky+�ɏ��>-Ame���%Z�Ϡ2�`sph�QÅ���[�@� ���G�װ����_���\*�g�-vf�3ыk=�3��ξ�i����u�9�1����9� ]�H��� ��cj'Zb�w�&�&��R,n�vw��J��x�#�CO�F���õ��:�t���� ?�K�F��9���);�s<�y�W�ft��>W�9Q��٢�s���*c���D&��̐a!	����^�h_���8Y�6%�:��M)jJ���b�n^f�/�{/���|��6��J}�j���eN��qq;�2J��|v�Q�
�R��R0��[�P�K��E�X���g�P$x�ca{�3�lh�#���g~r2�^�S7�L��CO�F=k�}*"�j�%���*@&��s�u�F��Vr%���,�cڽ鴇R�k0��oG�ӌϺ�&�,�G`�̕L �>��J���I����н �v�bX���em����I�t�q��K�G�$��݌0�~4)�i\�"���7�|�N+w~?�;g�fdL�L�It�K�x� *ޙ�!r��"������2��K{<K4ئ9�P�T�1
�̗����a��sO3��seM��F��]�:ipۡ�K���מ�<MȂ�:�:Qt��C>U�������"�:�o���EC��8���id�G�	O���v�M�V%��%,Z�������+�Y�%e�Μw/��}z��;��X��<�Ӱ����<����k������"�C� 1�Q���^16}�I;;�7x^7�Sgι�^S��0z}]f�'>���]q�0S�j��{Eą�=^W����� uW:�%e�u,�v���,��6	�Q��XJ<����a}�e���	(�TeI�)X�9��K� g*�9/�������y�Z����}���	 D�ٱC`�]�p��{_c���0y�*r�`���r�7�~ۥkt�B�+�
���o����e�	rJ\��a'hv��������@���r�Y�̏�X��B�Ea)+����B���>��\��j��\�'������yXd{&m6_g���)��I���ԋccg���t"*q��U��]���Z���͖�L�E�~��0!��v�zC��=,�"k��j��[[��3Þ'o�����0|��*��p���kL�bN���Lڏ��˳.J1P�A�id+[M1�x"�{���(#��d#e�>��sE� $��h�UXB箪ָ���\���I���`ї������'
� ��۬��1��#����^�z�jd��0�%������w�IA)n��0�z�<9��;	�F�D��|�D�a`6��:r��E ��0V5�0B�P�l��v�Ƶ��,��=.��3�59!5��I�8C�������JNۦf��UoֽD�}b!۠�9�r��,���O�vQ�����ocMD����4EO��o��h:	e�H�F].-���"ޡ��ޑ��av��ӱ�x��Y�&mķ���#�����~���_+�����������W���.۲B�C�'��d�*��װ؅$�^@�A�۴Q�L��(�j[B`�Y�Y��t��|��85[X��m��\]��w���YM�b���$��his�;�7T�_��H�pXbyg�T�k��I����PU��y�^쾃�`T�;L!j������DJ���BY1#7C�w���"2�?2��(�7 ��*�0�I0�󤅕i�,�?FY�\������*���s��1r#=ѭ���г�I����"�Qɉ�H���8��RY[�Օ�}3���7.�[�F:͘EE�+�I�[4�1��5p<kي$��,y���{�s�XO?$S!��}��RK֭w�ˏIt���jrH�\�榢܌w�ga����]U�T4���+�����J�V� ���Kͨ�aYVqԬ�|l�����s�'P5ք̞��@h �I�ju���_�����{��&|#�B��� �O�]ca��ϒ>�t9�O!J}�צ��|dCq\�K���8D-7�>�;3y�wyi�
���%��,��^,���o)H�	��t5i�Z�T��I?���c�ʁF�ܐu]� �,;�`=��+1� 	v�9i��3��	��c�b�S
���m���d�D����jh�
�;�~���e0}��)��~I����ϨBmU�����֎�"�'�{��nh��pMzPf��4������G�����Yw�j�-����)�';ɩb8Q|���E�`�&�F&�3/��@(;��r�O�JT�(@��6�?B�=1cʣ(�YC�X��&�榺\7�1Yl�M���/f�>J���T��N�t�Ič�/z`I�P��c��I��[�U7Q�)ace"��_�2y��� ����y����v�t@�T#X��Q�ѯAG!I�4T̹g�a*��%-v��m��L�V��� 4�Fi5�n�<֒��a��P0�d�WV���X�"��:
^��
��jqW٭Gc��t���28O�ײ�I���m9h�?d���/[� ���0��M���M�u"u�W��7�Ȕ?�������.� �<=�[��� <4@`����9��)k���R������Mq�d1�`�_�����
�5+>�j�[�\癍�^�Tp�����D�tN�xʦa���t����װ_���s��t�Z�MuT�&�z���0 *���s��|���4(l�1$�2}�/����c|�/�cz�̘�H���v��TE�|��~_��� �:�!O���ַG�U�=3�ke��y�"#�*d�*�,?@�6t�#�KM��@��$&AJp���E����r��Ӝ�z5�뉕���Ek�g#WB����g=M�̋��R]�ڻQs9�b�u���w�5��g�X�6��,8�A��us�I�f2v5-yh;o�#��D�K	�QL���d������M�ir�Hq����aOG�l�p�Jlذ�#M'���a��4��s�äزB���ogH��>2���c
T}��O�����OW�L��a����/EXHN�ga/�̆��Wo�m��ܴ���c�Y��S#ɵ�rYő���X"o��=�~����X�w~��'͓�Y1��>N�����m�␖�ۤ�,��.G^ej��,R�����T�ݓG�f���΢��\�0O�Cl\�T��/��k���pS5�n�ˡA�@�LـlӁ�W���`pMr!��q�X�k:Rr΀
��<�'�ǩ�-��h ��[S�U-�@1�����x��I|0 �/���btݾ��)b)w`���ZU:��o�&Y����6�k��]����=]0iF�a���s�F[E���Yb�P�E��j������o�ќ�VU�/����� �{��cH�0���vnt��ԗp�{xX�ol]h�/�~����|vt������W�ϭN���+t������HABWE.��;`�as&[WN���CU��gb�<ə��J�4�b7��刑�nx��Ҩ((��2��8"���]`%T%��T.Ù~�?Xu�U/�u)�F0��8���ߔ����J����j�)��6���h~�\�Nrn�Ȍ5�$f�(�ѕス��9��k��b+ڹi��sO6��V�lv��[:�y�.��N֟W0rqr�]F�3��'<doq�mPpS k}�db�ѵ��@����A{DgH=���{D$�	}+��G��e�S�l�L���'�u�)�����SN\�PE�/_��B����[!����U=%I��^��*|<��,�ϲ���r�0l6���ݕŨ�u��#O�6w`N��>W8�t�����m��E��r�E·����6�λ7Ec��5��\�����+�GfB��W���X`t@�����A~���<�޵�#$%YNk~-�}O��K�YE:�
��8@��*�ڎn���xw�e/���%(�)p���gl'�F��&�YV�Og� �0��6VN��7ƅ��
�!� U٣��v!E��D�֔�<c�SՖ�B��	RK�X#R	�N�庱���t����*�r�u]>��|���7۵a���;<P�
ޗ>[/)&+�4�s��A����Ӡ�Q�R#�~�b��6!v.RiIC�h������������	r�Sy��skM�#�f O��SB)�	g9M�`=���bbA�R�w+�<�0`Gd���Ĭ�s~t�&)f�[::�\_�[)$�9���~!�P����Om�qSg8�����?����$��B�?Tݡ��N�l
������5���N�1f.ǲ`�d��:�64P����Ye�U���/�Բ�{���S7��ߠ�z��v4D�9$�_V�l���i���璲<����J*vI[������Ӽ&�#��p��1�fv〙4��f�vk���7�Ҍ��w~�M1�خ&s�r���^�{���3�����`x<�b9���J�q�M"���0�|�:�=����0F���v���p���+h]{��`$��hO�|�.م�tg��P.o�؎$y�ފ�60��{�6���Ŏ4��L�����NOǤ�5���K�Jԙ,��=�I���Z]��%�UC�T�/�~ڠ��vI���j�jDn��2߶��pN{t~���X�߀w\5O�S���.����_V�Z�!0���ꕚk��g��P�/{�|r��>�����(�2�߀O"7��N;�Џ�Fmxd7�a�v�����P�
]b�M�=9	X~:e#����-�$���po��~_Mgyf�Ŗ�W5��ue�LJ�R$B�U5i=��*#��[6Z��U�>T�#n��n�EPdf�?n�i�$�E�{�Ng�u]�Bf�
�,�Ĉ�(�J��lJ?Gr`C��Vm'�0��~��m�݈��4G� 1o�1�{����H!���Y��B�Y/����<u d���1��� )��p+��7�+M�z�7�C;�r����G{(^c�[,�؊��XZ��s��K�EK^R���^66)%%�Y[�������n���c2g��(��.'e�&}t���N�W���z�v�B����;�O�[���2']�q���h�_��?�Q�{�M����S����SB��l����&�9.��ّ6e��D�+T��0�c+���c�PF@"7Y�P�W�/(�`��S5HNT��k���˺��3�����t��fu"4��t��]�=9�%�h3$Rt�Dg������A'ǳu�4w��l4����V0�̾s|�X� �{x����"Hا�?KIb��({�����#|�f����Nl�O5*f`?��<�:Mb-\���a P��ޚ��}{�X8�"Q�<F�������կ�]�P��=0��v�oy�&5����%�<.���'�p��!t�umx���-DX�����a�s�gJ{���T)�Zó���)���gH?7��"�"�j]s��D]�Ԋ?��%��Ȅī�����E����6����!;��/a�mw%g;	*�I<�*TE��e!<J�p�|H��Y�qW��%e]>k�˨Щ�ѴH�/KZͷ�mF�@���鑉,J<���[֢�֘�f%;څ6]�yx�7�����0%'�t��&} Q�)3�K.Z��V*��-Y�wG���҃{�dS���@�x���n-��B��+��+[t���ڃsn�+-� jh�ܵ��/g�x���>*s��� yW����dm��۷��<�Oiy� y�a�Ĕ{�/L��y<y��e��+�v>K�Dܛ|:�1O������lV���k��~͵�m�3;�]�@� �[;�qǎ2*�XA���&�p�;E�ZX���Mp�w�󓳻��>��-���ɚ3�sG���_�@�����HiJR�I�C�m��@��!�Z���I����3}x���ؠ�|+���r	�EQ�H�S߭e�x�r�Y��ܞ޲��+of���{-|~KG�u��?���\�nō��AX|�g�Śi��*0%n��˟��.��m �B�W�oSC��OJ�"W��Bh�x�3E*�e�i��2a�T$&i{i������ �y�}Ҭ�&}}��{1���9���v�g񆌆-J^��|��LN���Ɛ�~������W}D�k�TrT@��{3�>��&ȥR6�4 �&��Y�R-IF�
�j�ƚ9�#ڻI��F�h�0a!��6�/lq�-�X�����Pwn�]��_TV,�ц�E�J���_�Z��z`*���ј�b�dqqk�����E�*�~^���ǈ���ERu!�SݛN�������5l��V�׽��/ho$O]ii�V�;D���E�?ѿi-Q����E����-�>��I���z�wHDǷ��O�
��lEC<"v�%��F'-�C��ѮUJ�f���5)���4ݱA�dFL�F�#(�7��V0������c��P^#���Tb�!B���BS�,T�f���}�ԗ99�O����D����[�t\A2䫨����[D��pb�':���M�τ�}_f�ňc?�R·���5*�ٹ@����x+VML8��#��Ğ�[�mJ�Y(=3��2/��
$�MO8�;���2ot��n�1���'�fz/��Pn�qH>�OM�~��������������7T&�5���a��Z�{���ԋH0�����ޖ�����v5~gת�^\�.ɤ�ܠ XT	߷ɟQ����'N�k���4�3V��^5`�ܘ�v����"�Qt�i|���{f�PV�"��xW�.4::eaݡ9���ĺ���@���k'K6��9��~������+���\��tmvI��9B�U+�5P�VB����$��q��,����խ��{&Є|��E�24�P���Og~}0Gl���M�ݵ��y���C��¡�Ӊ�t�����Y�s
�,���lx�fߔ�B��&Cg���W�rnD���7K����5j���)G�� P��w6^ \��5�wU$�\'.�-+�\`�l��X�\B-�1�k,��6��l�	�5��o~.BB�<g������&�q�x��}G~ާ�@��rr���9p���rq3��{�Z|���n�x�5X�#i��<Q�3�^冪������T9���u����!xhm*��|���� ��@���~�T�F^��;c�k�f�C4sr��f��5����q@�K�����ð+�N��9��c0!��'z 2vG�+}>t��l;E箧�W�0ysM�&+9{�	�����Й�0c��b���4{<���
��y1焟��;
�ۙ�=�̷]
�?�y��thD;�@s��⒎0�(����cZ���PV>�N����^�Eߗ��X���d�pP�	BU%��-�a#��;Eɼ'/��X��,�f�ѧc�>
Z��]@�����!GՎ�U@�Ò���")kS��]�q0Z�1��OJſo�.*��h^؊��C�:��?�ڴy�)3���BPB��\����m��Eoz1B�VpZ�tF$�
�3�����ǟ���O\mv��q�)5���4~%�@�DG�1� ^n���L�-�1�Oc��ŝ~��}��0��-��ôŗ`��z!' �"mU+��>��Zr��ʿ|C�tߢ��s��hs��.@�7��
�aO������ҟ�+�#\��F+҆�.��}=�i����2,F���7�i��W�S�MJ-og�3J�U���ںΒ�&{��Z�Ɇ�� <ux��® Q�*���ޘ�5y���Y<�X�1����9)/�Ԅ���8y.�=0���7�3l��zR��0僆�l�;�Gx����j����W+�� ��k��߁-�QA���ņIy )/������i���>�r/+��a���^��*�%&�Ư��$�$D���Y�iS(|�Z1�x���"]#�#�f!�V���^�Pb���B�`dn�'t���L�r4��?wxs[�A���*����!#
B̛{���*bY�u�v)���ɏp�":3/��-�����5<�jR�7����<��[�m�77�����P>)X��Q�YVQ��֐�y+�CNѹ���fG�@�d	SR��qc��kc��[�R��M�ﮉͼ�[���H�Z}�H�!Ѵ(�y���븨��Ԓ�˖d�q#*����|nP�,�%p��4���J�A��,<�u��D�����Y���Lmu�`&N#Р�ċ"aʛ�?����]�xP��i-`sIM5-e���;0��n=#D�$�Ⱦ��:S�%,��jL���I˹XK�o�����1�|�{Ǉ�ҍ�/���8koyb�iL�[�rm�>��d�JE�N{�|D��/����0���HM_�-�$%� �Y�0�������q��VoUI�?���}v&{�9�t�wȜ}�2CD���.m�"�6��\iz���!�a��ȲuS�p)�������L�v�W��chq[��ѺJ	�]a��"߄J7���o�h�1p�	&r���W�m�M�,���*�ݧ�C[�9ߴ*	��[�wE�:�������D�/@W���<_��ʹk/�΃�ݏ,���#]�t�dPZc��B��S�]7&����o �� �ȧk嚌ر���!ڿ���7��_�ڙu�����$>��'BR� ���Р����7��F��).���� ��h'ü�f02�4�`j���Ҁѽd�'3�\�FW$M~*���V�g֖\f�����'w�k�p�_����:@$��<}[>{cIx#{���&H�*c��^R����s����?��  )��p�}�cq��
�DIøZL�^�+�Ϊ�����i��*�KL� ߭={���?���;��E���K0��$�
k���š�aPj{�%�j��m-�����>����b�bm���m@p���2�Lh鈤6��@��B�MqN�4��O�Gv�r�>3�'ZP���]^�K�| %;��k�leXR���5~��*y�ܳ�� 1m�b8&�&A_M�{��$���;$�X}�y�a.j4<;,U��\E�cx��d�I��^S�f֛��� s]揗UA��PI�<��(pOF�{q��e�R�qG����ś�>;�ZcǷ+#Dg���C��@�sٸn�n�n���F�2�.EL�>�?�o���tcCy��]-�t ε'���t�]x%���r�g��3����Nt9�a�EB�m���qt��h*���llL�Q�����I���	�r2�:����?Y�*A�����{{�$�Wm��TW��=bO,�	L�0q�$v���9�yX�z�Xı9��+�6Y$��5�C�t��W�sɿ��f�'kA`0	���!x�E��mmr[���2G��=
Q�+״�42�h1X��kb��1����&L`ri�"�UdɅZ�4>��8�{�\E��pC�=�zMaF0��;L�C����WW��-�y`5��Y=h���P���<e��fN��L8��G��mYl$�_E'+����%��E����`op�g��0Ў�N���b5�N���8��-��\Zu���,|L�/å���5�ɯ.�YuO'o1V(�:Sř����9ty������V�y��%�,86,֞E��ڞU��D.���h�}�6m�����ɓy��6TLbet~Zq ��r�S3�L�U< `V��� ���ʂ��Hth=�����41���%�=1�_��v�ɼ'A��,� ���P"W
�-f�+K*�!�d�j�a$�8PĿ*�}ů�76����͇�ٔ�������tk���4�z�"�M��L���?��~���{]���7d��v]:��pŔ�A�Ago�I���C��fy�W�&;'�=/#�L7���^Rg��}��U5}��N�] SC1�czOߍքC�46����S���DI���d�Ej��]X#uvL�e}SF�P�o�f�� �('���Ū1�Ó�?"�U���0^����LGT����)?�"k�EU޳U��*pt���U�Wݵ��X#b\��A�17捳�`HL���!�N��`C�Fq�Ev>��1w�7�Ki�g��4&���V4�$2W��������� �Ll����ڭp*.��G6m�z�G-��u�*�q�\���\Vy
��1���<12Q:�.V��\�����%�F�����-���=�G���٬>�E=I�1��É�K�\�ʹ���ܦ����Ui����3��d;������'t���ֱe�JG���@�bCQ��d���)KE� LZGS�*(�O��o�3fu������+��,����<d����{��=�Mᮛ��(�4�ScƢ6"c�hi
� ��׬�{�`u۰���9q�������9U�� e<I����a����.�|�WMԮ�g";1�µ�f�zaK�z��B�����I?c�o��q�Ʊ�H,���6_ |�ox���kzb���`�D��I�Ԉ��>� $h�87U�;�4���{T�̏�#ј��.���K�I �`��Uؓ8	���Џ@�u&4h��Y����]H��(�4��	Xa��]��v��.�
����Wu����|X\K� ���uP���=����V����"�V�t<�B}�Z%?���7:��X����B�ڠ-��l���N�h4F������ԁ1-B�)g�y3^�A�dF�����jחa��(!&35�Q������o���P� 8����&-U��E�Jk��A�<��G^�>l=Ԟ0ΕMۑh����-�y��-�he���3���٭�$�_r���B��27X���њ�<T�I�i(�)[�z�I��=�<�����Kؐ�y|�l��=a�m�_��j���l�����9�݋��)��m�l�X�>�!��%!���84Jzw�y�*�Zo�1���%��'S3�y���;f6����4�k�7�͇5�՝��2
��\����7+�}n�h.�	]3
�b.��R�[Ҋ��j�M��>��i�A���ǟ$_ɞ=�_Q�,藂!�7�
�ne=�]�h��x`ݳ�%fj�Vp-�7Wq��Q�2��<�ӮFI�sm�&t9m���J���
��wwk�3��bMs��b���c*X�4"ߪ��2��.(����;��>+��S`��s����BxR�a��@^�+Xb���4���JHR.��� �W�����}^���Z���R����6���ղd�Ń���:�O����;��z|����Z^w��������{}��dtg�96�1a��ȑ0�D��� 60qU��l�_E��&��^H-�dAn�T�	�T@��nrP&���gۥ�X8�i��T���:�@��y]�~����x_��� a��J/��%۞��b>Z�)�"Bj��G/sF�=4�螑�V��+���[^�.\�?����GT��=���!Ƙ<��|�V����c�<g����빞�@'O�
*�/ik\���8?�m�>9��̈́�=�O�/JB����8�s���F9�H�`��ţEFǞ(�6 ��y\���_b��XJ'8����c	���<��7�Nh^}V�ZEy-�]�|.�O�t�ᗹVO��
�,���%0��v��>��w���'�m̱�����Q�1q�Z�PT;'y�Ch�i�{7s\�$�	ݞ���u��M�Kd�$���?`Z8��U���Ѿ���W�7�Hz�� Yk��Q�(�>��^���y���LfWrf�k�����9'*��NTT���_�� 
�J,ഷ`u�L���D\���)t6�wk#�bh���ʅ�&Rʯg����^��?2-7����R���'�&>�E��7�'�v��9����N��.v�MRyT>�����{�� E��˼��p�g:1��H��N��������cA$���Q9�
D�7�Hc�}����}j�;����B4�Ug14����������.y��rG�EA6���+ap�ZM�먆����1g�Q���X}�~�sk��u �O�Ձ�(����v�!���G^=6 �?"�-.�M-���8�+�|4�v$�)e�z�6��)?�p�X�p���cU�D�?e&%�[*MG]����fP�U�=��t^��]q���q��b���خ�����c �o3�I�Bވ4��� ��֕��5a�R�M���A㕹�c�l&�TZ(�v��u&�ɫ�+SG��#��:\���"��"F7����Q�o�S0��8��:�\�7��>�����:��e~�:*��j`�e�W1y��S n��;M��eE�2��Ŝ*����Z��4i�h�SH��u����Y�����"�5���8���@��b����I�VaLn�?S����n�kn��> �F���U1��:K��K�n��YOb\pl�2p`f1S�:�Eo<3�E����@��A��y�l�J�h�
���/�5�b)�4/���kdd�5\�M���h\+G׺7���*��\M��L�rJ�U�oИ�p:��'�ao~�{�Z�"�5[�3l2gЗ���A~���	yv�}�V�;V1�H�[�DD|L��;$_��\hGX+�kl��/�LI��tL���0&6ȯ�3��#�I�s�}r��9=0��o��^�f�b�S��T�b�e�}Wp�	���P���o��4yX�xC�[���b�D^&u�H���?�ټ�CAӖu����"*bcV��Jgv�d���C	�n���~֐I��o �����Dh�@F��5�0(�Ĭ�Y�v�֏�Tw����g� �Hd�p�/��c鮺��	Frr�ë!s-[���{34i���O^fN�&�l��X���܎���&^N�c�ű�����,v��!B�3lg G�۵���FN	yps�4��,�9z4N���c���s@}���B��tV��du�y��\����ʾ���a��@�^&o��\�c��"�A_\)�,Ԉ!3L��	]�1R�-�������^~�A�<�έt�����͆B�q���v�P�1�5T�hz�$������TtS�ى4���kh�(,����Nw����==:I�^Vd�D�d�f��0d�ɥa:�sR��+Y���!M<���r�b����Ba�DD����գ����Vv�6<�� ��_��ĝ�\=��y�nA��17
�Џ����KP��пv}�9H�̕<�|��?{ ��.e��I��[Kq�6o7��eP/+l�a|�e܅50��x2X�1�������W-eմx�:yDF���9��Y�������Y_�W~�O6���9.�����x�bd)�M�>��3��O{*(�ƚ&C2fgiS�z�'w��,��c֙Lfu@����B@��Ob�ۙ��ޙ���g�O�S��Q��o�+>���.�)(@�������O_Q���V��#�(�� 4�v4�r���w0t�ٲ�[�.=���e�s�#��/���3����� �������N��@ ̏��kh)�?�<kɢ)�������+1o���7
fsX"�PٓYB"�>7��U\͒��R��;`���i���l�ő������nQ �L2kR|�(���.��wfN��h��vP���(��GH��	����������5+c?����Ӆ�b�p������#�!7e��b�?��^�A>x6p{\$�vE| �'�3�����?Ow��]���5O�^&���Odv����5��������!���� �pލ3�"�k�z��u)�}�8��7�T*L� �) r��sc�!����Ώ_��p�#(d�aUpp���7@��]�%y@u��-h�>@+!�K�:�^�(�H4Qa�����H�]+�1�8��rⷭ ����׀0�\����b#H�Sʣ����OF���R}��b�g�B2�� �-ٽy��h�؞�ɘ��bs ��J-h��9��K*˚�Q��^BG���{8.��,����Gʶ�T���@?.~�y����sw��A�b�x�$_���Uû`�J�#�@�������3+���\�*�e<R�	��?q)�l.��!�i�/ۣ��M��ښ.>[��mM�&�LzC�J��*"�����1o���&#�{ɏ^��V��ճw�� ��F�lJp~��������,h�naЕv�~��P#�1!K���ĝR>���
��Z�\N�h��[�6U�����e��=�����(%��E�|���9������
Yib�*��n?���G~���;y1�W�J�1�w�*k��Y�M�g��� {�:�>2�)9O
H�d�Hv<�#m�B���<���"qI�O��W]wF1E��<�]�Y�bT����0�%�W��i�bn�Jh�^4V,�+n}&u^Ĵܨ5v����*�cq�V��BStU!� l�4ˮ-��Y�}Y�턪��>�-g�K{���|�KU��g%w�~iU6�2%�0�����O�4rp0��
��������$͡iN]��БLF�S<s���KwR��,�ԅ�.!��1�'Q���k�1�Х[�ظOP���	p�Ń���H=ʻ0������Յ��I����A]Cߦ�|oi���z<�mj�A�%3����T�G���"�s5�4�t
_�C��%: R[��/��U��;0J����h�`JAH�z;���Y)�BD`��P�0:Y��̃˃ȯ�r�y��e�R�G&�� }Dhs��N�z�"s��8X|��l�|9�4�^o�^�O"3(7b���'��㴊�ܦD��0;�֌9+��[�l7�0��%�	]�%�)���K�"7��]��oI� *�1�il��i�@��:�k�=C3!b��_�NlKN�X51��[o�4o�ld����/#�-=؃D3J�~�$�׉B�ι���{�g��pRV#�C�@�^,��V���`v�(c0�� f���ʟ���N����*;̾���	��'�V|���������g�-��"-�.^��&Ov.�x>�47��C��:!o���b��ٻ�>�u����{��a��;��긟��A�Qy�Y���õ���Rz��J���Ǎ�I���n���؀������P���_����?U�����b��T�Vڻ���qBۍ�?����1+���nf��ǲ�Q�3膗Y���@�`��V����sF�w�RV��ߪo!��I�R	zQ��d�x�w�lSK�V����ּ���X�-dï+xMNIQH��r�6b�gkm�9���i�4_�iK^:
VS�ִO�d����w���������d������9�蚞�T�TcSd	'$ 5��d)�e��ޅ�CBBr+Ҕ�K��Oi�isEA��ǓD7Sr���8Ӗ�����3�)��9��s�<^�I�R�����-�q����z�Y$��E��[,^?�mݾ㛝���{�ŝ���>��v"�ۗ �x�I�OvtZ�y >�{�y�n�=��:��F@�R#�>���Р*n.��!��*������wHO�u#P��/�>�^w�g��c���,!J��_)9�w�%��Ʋtׁ�yp����`Xg�cە�Â�s�t�(" �x�(e|9M�U>�_���r����U/��hX����HG�ᡦ�M�޾&�;S���'z���E�2K�q#���0Z�T|}>�1�[��<l~,U���ů"���Aѷ�*@K�m}ٗ�۾I�]|c5:���F�7�:��,����.�c�_�h^������y «�!_����֦&�}BU2L�`�5�QK��I0LX��D'�t*��%�8�� RF�������P1��GĎs+�9p�(��~T
*zs9�;�����8\l��f�X�s�.'V���Zju����UIPD9ſ�ō�ժ"�oS�d����|��)Z�Z ��)�P��C�W!�g�xR ��S��J����/�]a:۟W�B�VxH7�������ke�o����{���N���_S�`�eF�,a�L��4�#�6W�2�	�>f�Ԃ�W�W����L3b�/G`!C��h��9"���.��	��7�su���Bd�I]sQ�PN��Y@�G�O�g;,0��~ş���$;���N�;�č�h��ҋĚH�E�A��@E�a�!_��J�=r�iJ���A�I�8Zȩ��i�釁gC0Ŷg~��%�*V�A�c/6SX�Ԛ�$�AB�x5e=Oa��x��.�_;m��@��m6��hI�/g�]�M�s.{ЈH^�Z	�jׯ���?MN�� ���S~���� ��.�j��ߙ1�"S���
.��Ҭ�l �����$���3y�N���)�ҫc����.��\,�O�c�x��v�\)r��A	g{<6U��ר-�!_�!�sN��'7{���(�9�Cm���A�	[���6{3���l�d��1TS�o�kyN�B�M��*���޺���D����̭e��0��/��ծB��a��� ���,S��wX���:i�����)���bb־�f�q�w�u'�+��gV_ R���gO�	VC���<����v��R3��+�m��D��-��ni���)~7��k�Y>V����Dm�8����H�*�Ό�����_��7O;��NlO��nuq
n~��qp�m���C�N�8�����e���b���~�����(������V�e�G��4>�W��Q�V�+g ����P@�z�HŦ�n�X�3@LC�m�?�	B��9����Oda��)�(�`O��%ܫ���
�h;�,�о�Q�B��u�X��-^*���])�8n>e~�6��!�p���;?�g�M�>�9k���՜c�2�[v:^�
��ud�`+-o�����ծ��fg�q�_��(��S����kK5b(=�t��9�K"p��\�?�r����θ2�Q�@�8D���|��{�Ƙ�kF���.s��j�?�Mo#^����e�(|�s�Q3!���H�2��Л�Q�/�~���T��%�$�AP�+��Fl�
Y�e��L/ d(}�Y玺���Qԃ��:�N�h�%��4n����x�B�'(J��?n�Ԩ\!���w?�яzk�K�r��jF�v@h�F�p	�?r[siL�2sx���xh�����_�q#f�1f.��?�m��ݧm�E�PZĠ� �,D��������o2k_��K=��<z�>/K�Ue<��|����.����>.���Bf�?�?z%}[ �ע�L`�Q�*گ���X��<Ln!���������-����T��^�7�� 4�٬�{�R��vݒa���WKN�fI`����(���lbɞ���\X����$���_T���jh"�etǵ"�f�$:
������M������'��J�Ħ�4�����K��~i�P��W|��%e?���=�A1),.�c�l���8^�%�Ǳ�?�IH�;����9�;v��n����>c,"�$<�#������s� ͠�Ѧ�DPo,�m`�osݳ��<�e�`��WP0ӳm��:�I�%&JW<��]�
8xp�YQ8?��D��6��<�k6)j|��lj�	/����55|_o����Vi�� �N��'�5Y�Ŭ�"&�VQ�&BL\�#>1!+Tp_� �GN�ą��W����cf	.�@�ermA���e��}�>"�b ���,%F�=�7���E�;�_����4K2�V1�f�]����3Ѭ��x��Y(�E'��s$�#�\ �]"ۜ6*�3�Z�f0�Hx!I�VmmzϾ�������W:��4Xs���E�&1��fC�����6��ж�W|��i	�-��#�0{j�ѐ����}��	��3l|�a��ʸ��3�Y��9�a�辋�G:����
_l�9i/��^.'ތ��kz�|�~P*�C�d��+���Z���(��/���l���HV����g|���(I'8|j���q<�['�9o�jop$���r�U�����k�$���.�mE6ĲNG���Qad-j�'"M
�[q�aV�Y`Bs)���q�F�H�⩡݅~|��ʲ��6'����I0�k;��n�b"��O�h�Yf�!�r����	f]
'�����tu��v�����5[ZN,s����܉��g�Ȩ�d2pI�#cQw8j�p�:�y�+6p>!���t@�qy1k^�� g�[A���@��w)�
�c@B�U�D���6����L���G��4�[����:~=�C��U�;��>|�!�W������>�lN�b�.kP%0�v��� ���_9���{�W�)�گ�O�Բl�������� �mx�唰�1��]�;\VV�z��NiR��;��J�M��gz$}����]��܍�QT���� ��3Us�H��*�"J�H1ތr�-���ո���uJq$�.#ҜT����\+1����'�24.��

������g�}Z���,`ӄ���#ɣ��6:&��h&:"�٨N=�;�*) z�,����
*����#����=�&Q�T^���D�ٌ!��U�$Z44�׆��"��б��a�]����l���r�biY2�P�ofD@F���N�x/A�X� ��e��<oL�ǮO�;^�{i�A�?�9T��b�������Q�t�����m�t� �3}�Pe����c�i���Dpݖ��3p�
8W6fCw��+�3BX#�_��5m��y��z�v��9j�Z�e!�3�fG�n��'(��Y6(w�_h�Y�p d?�`m샸�6 u�>5�����G��#�_*�<��b�V1�*w�L�������x?���'^|d���ѻ��F�h��FHUu���o�+��˪V3���;�"��hu����Y�ݙl��0�tʅ�+�NW���e�G{T)��?�V��k�J�p��#��A\o��s������<��A��Τhh��AV8���m���n���q����� B������;-��9���OVm#����o��~VB��cyx��mU�5�Jkc�\s GЈ//5'�Y�2���\(p%�P~�'��d^�f��[��^�a*��.�2�ባ`�0��H"�yU�\;uDl�Y{ݛ���wm�B�p.P�@�;�2���\��5�\�J�	�ן&�V�����9�G���#��[�~��Ј	�;��p�Y��%@d&��j�3@��������!kg����4�������pp�	�B�9-��Z:��qik�|�%m:���yaU�L�
L��j�3G.��gO���O�S���av�Z�V&l����Z�]o��}t�bi��'v�>��W_��O�s��t�7�i}����-@�v���2��dA��B�N�Ĳ��:��D��	-�Qj<p�\i7�n�p�˅v�p�u ��a�X_�!>�^�����-.�� �GBZ��������^���[�2����i�6(�*�Y��(^���i�������ϔ���qn��(��������Ժ�?Ij��?Wp[T<hU��j�=(�ρ���D�pF��ܢ6O���O�����̝cc�D��xY�G/x��j$���p����/EG��|^K�������53��ź5#Z����4o�ߺ=3T��G��FS�W�(:��\��כw��Sl4�l�&�g��W���B= ,��|��y���#����];�fZr�u���l�o��mD�+�g�"OԼ���A?��U�p�y�������/l�)H�YF�Q�`��`<�!u���#�s���K��g�l�>瞮�TIA��Ő�U�E���(��'$  A�����r�-"/9Iً��&��i��p-���]��?t�؍+S@�"hOD{Vs��s5v�$��9�eL�2�h��h�����q�?�E��Tk=AQKo�3�y!��t��v}CU=WG�ce+#o�gU�����(�Ź�Uzr�]S�!����Kӆ{�`P��
p���~���,���`H��������Rү��� +�[}J0ۡ��e�>�P�3�OA�rx�6�'�Yeg-kJ�>�w��{���O�j�d�\��$APW�k�]hZ3s\��� w��]S+N�^G��;�d�I�M���l� h��լ�Ax��e��v}X!�P����P.-0� �Mda�i?4�Br����� '�Gݓ��ݨ�Z��	�e6�əQf�#����ᮍU+˴v�,e?j��B�%�a6�BE<[&�[{Q��1�pކp�'!l1�J�Qlw�w���g3��0�y�&��qZ����݅ �|L&���1��af$=ƾ�If��|V)p�6��鬤�V�c�$P�Ŧ��KT�ꔒ���H��P8�W5�?�R[��F̴�LD�j%�(�\�ZW��.�;���Q)(�f2���_����Ѩ�d����P]@�7F��d,&.���5�v�n��������@��i������E|�(�����c��ΨʀHy���wR�#�� j�)w��I3�����lt|'x�����Df:,@��W�B��e�ر�P���5������3Fy"��Ao�b�.D�1��g�,6+����C[�0���V�[��1O�,Lvy�a��3q�vy�v���O׋�_�ZbKS�~��vz�;]��GQ�Y�i���)���g$R�k||���Z#�C8�����2���3��27�҅�S8�K����������zdBW֮�5�T��&)�\�ny�Qy;�BX|�I��jΧ�4���֌�W"}�Ϊ0�ءb�-)��KaVn�3�>7K���Uz4��7��ݐ��V��گ�Zh�]��$#�����x���DOQ���E�aaR`�6��Wi^Y'�B	���5�ݐz�������7���*c���v�]�	7�T�q��jlBxR��ԩ>֦��Z(�R��)�{(�3]Im����;\[�ӮZ�ź*���Ft?�ݼU�֮?<ks�4�I>�%�s���Yė	/�E��Q�h�`u�Ǵ�a��$�,�""�Ě����X�1�a�;�ɜN6t�<��-�9İ����D�.|��������Vt�j�I������jF�x��B��WԤ6�
5D���$A�-�F��x��0^�/�8e�B#��=��=�8=��ƬС���(,m$#�l\�wQ����>�s���.>`eI����l�fζ-��J�;=Y���9&��Bi�G�W^j�D����8�)�"�V�or:��Zw��F�]=�;�׍*%~�M;q��I���Gl�c��߸���(��PK���q������$�y�Ջ�+r��h &
��&�#�)B:�,���bi���Z5cٔD"8�+V0����ꃴȲ,|	�����. �*�6��-T�5H�]\�2
�L[��rC�b7�^�?�IV�lƆ�e}��duؘ���K4�O�x���f+O3�lcP�� "����:��w��` �#.�����
���e�W��)�1�0�'�E��\����Ja�,L�� ڽLAT��wF㢤@�$5Vn�0l��w���i�`��aa��ګ5�.��������o��Qnn����G��l�\��Z���A�,��������{#JY��CC��o��D�og,�-�#��8>i�U���y,��գ�)3��@�)]BbK(1@�@(p*aL��A
01(��q�,�Z��+���8��xnr���<��\7
�y��-	|~>��f�c~"ǣ�<	;ͳFE�e8����&�j�BPR�4J=n3�ޚ�}V?U�T>7Ź�.0�qi|����A��ҙ��2^0�];�EQ�P����'X����b���j�:��C�'��ͯ�:s��Q�y�D������d��(`^~���� �?O+��A���6��Prl�aʔ�~O#�	k�\�Yk�ȚXCS_�2�ױ,���Fڥ�*٘2�����_)���BK��<Ԡ��u/a����E��n�� ٨��V��[^i�#�	Qy�gv�Upx\Ra�/gy�Y�${����`���F�y1���$H�_F�u��n�&�-��ǩ���L�<�R�a�o9N��+ruQ�s��q�d�.		VVqb��R���i�������K��dA�:��&�G���m��U3�3�����Fo����,��� �w"g>����r'��»�U��'`5�r�d6rEm���;/�Y���k76Ͼ��7nn��<Q�i�zYۊ���k.�Z V&��^�ܡ`QS�i��c�9L~���Z6��]���h�O��+J4�3����
�,m����?�q��=ߔ�,��Es�����)ebe|����+c�C��w�*"<uAo=Lܹ?�.
�?��U9�2�r�D��_H�S�� ���'KȂ?���(�Ͱ�v-���a�k�X�C���T���r���q�]��'/%�*�8���N8՚��"�a:B.����=7W��yZ*m0(ג�x�'���2�_wĄt��үuS/��l�N��]�����"�ְ�[k��We��S~�K�G�t�Bj��p�i��<��K�H�I�Rj����yyG��n��1S�e�]���輝��iȟ���b��b��x2$����A5��O�11�BtX�R�;KC]�amA#��)�5�8,��H��7����͔�Ƭ���˰�%����b�~]���_�Ǿ�\C`�ϡŝ�VF�Q�J�O>����z�ǥ�kjm�Sx�S�H�i�����e��|ʙ��d����Ӻ1���	`��@x���m�:�*Q�}�ʒ�g�n�WPF���!�9���*��}mT$z��LGۿBB��d���؀�弎˩9R�!�*��<��j�9r���O�K�--���r��eA;e��ht�Fu��C��¬+�h�_�����=�;���D��2t"�v���N����aL�$FIV�J�[���C���a=
�ޠhX��G�N6��j)n87p���/1��V"/��)i�5>nu�,��,����48ό���1�\C	��5�E�Ԫ���2��H$2��H����y���۴�l��dfk�|��R�M�����B��+�����p6�y�+J��7h�*�b�I*r8����l���X��Ki���ʲ�� �93 #������mZ�ظ�����=y"@���d�5i7 1^R�bM�y�ytm���6(��|5Pz�<,�����TrI�υ=h��v	��C�i�J�_N����W���Ub�{�' G��4�4����1�I 遉�t�?�N��V0�����B�����v+Ȱk%te��o\�sc��Y2S�D0ձ�n�叏gz�c�/N�$�D4}T��.v�c���V7��l�$\#|1Wu�/���D�H	� �榎���/8�d�����Y�<ƿ�~8��cz27i�y�V.1�pM%�}M0�k��'�#W���W��5SE�I�6�0j��z����_���NW�m�`�1E�i�擟 � ���`Ɵ&Q��0s`�(z{|2�~�?��+�m��S�7�
�������(@:�~ϭ�coo���.|�M\�n�;v�����o��c(\2F��J5~'��aZ�����r?�%	�����	Tgs�\[�q����H|��~`�y
?#��T�#
K/�#zZ5�ȳ5�mq��\�3r����)�No�|��g<}���R�����9�� +�Y�1� �=D+4������U������/Lػ�UQs䱶8�Y�c�����.n�7��*Ƌxh��a&wB.�:#H1�cU{��}I�09e_���SH�]�gwS�OD)K`���W�]S��o���w�,t`Ѯ'we-��@K�0�?�~+�������}'Q{��z�|܏��{�u*J��,�bō���nG�+�v^�2��Q`9W���KH.�W����8��o⮾���+%TD�6�Q�_J������G}Á���Nv��T��������H��l�Tp�z�j�C���U�]��Μ�4��C:U+G�S�*<ja�m�zQ�{������@�s�_e:*����F��O�mt\�&�܎s��|0wDn�o�b�O�*���}�@x׍i_�EҨVLjs�^�T7��-Yu�O�Ֆ�o֣T���mht�H��p�#m�S�4�]�$��'~���zƛG���Z���������"a���E���T���9�Fd�{u�">���ކ��UÓfP/�lL?M���&	�m����)�z����)�&�ժ �����jB�Iѫ��D#��$4X�[��I���B��c�nb�S�P7 ��#�H1�]t��_��9�笻�C��\���Zh���[դ,�K,-��9�^M.��5Ǵ�oPj58>�Q���b��5�G"L�YC`v�[]h��)�~ahܜ��1-=5��̊&�Ր@ 1���W#��#LH�F`y�E�c���_Nl������+�I�1&`sg�Tp�W4�>�W���p�[ޢ����g�hفeHү.ϐ�����#��o��e�)0 �� 
W��'�;�	�%�ʑ}�������獆�ʂ��4 n�_�zPbߓ,=��_��p�|բ�C{����*��&/6	�ypO�8��F��R���I�؍�\�*s�+t���2���:��~�6���M�����=*_���B'��?����� ��@�L��L�}��J+���*�}�:�{YW���a9�|"_�1pӫEY�˾�.��OޕacO�t��<�7��j�B�����.��E]'��ti/�X7�����z)©���z����Wh�[��>���)(��D�h�c�(1w�ձ���
|�:N����y)�1t?�t#I)j��  y�29�CjQw�'4^��1�?:Y�i��X&����;~��[m�~�������Fĩ����o.>"�{Z�BS�uA·%�2�}e�}vOYӌ�#Hi���2�2�q\��F�2��D!���+��*��*�^���P�/�$��;�`�3���r#�tǺ�g.i+�x6�Ȑ��7ۄ:�IR0P��|u��~���N���|Z��4J�%��]E�[�J�ʷA�
PuW�#����1�����e�/;9IBϐ�J�]v,&�I���K��q��O���&� ��6�f	��Њ3�/j0��I�������͐xY��b�K�����^vQ�����ɇu*�P��F4j)~�!�buS�Pp���a����7=��"63(�O��j�`p��c�qJ,��9�ۢ�������QN��8�5�#C�-��#
����2A7�V.��E�E!x��V���bB��%L-�͜Ho�&����a%>����u"�DvN���$X��y��U^�$�Y��^���N�.�5z� ��x�C�D�W���Ȱh�M������:�|s�i�&��/ ^���lmM�X0��ɣ��dGxf鰮�s�)3�|ժ��	}
K�F�+/tǼ��p��{�t.�5�b�r�������Z7ߓ�<,<}Sg]���A�7B	�\L��������7n���T�3q�^��d<�	0��h(�!��&��x�ޗ��5�*R9��l�ҍ��EHK���̱��	�PI�%�`���l�N�5*���95t5:�O�����S!!I>��-J�&�|��p�4�dT��
��LZ��+a���P�c�D#rs��G�;Qí6��C�P�L$v�je�/E!���~}�!�Q�[|���
�� �VJPM��l�xw���ʦ����&��%:��Y�P�#��LDn�5 �|�ð�lE�aY*���ա9������&�k�^~�!�<X���/�m%��� 
?�:��㚗%}���gr��L#�=xƘ��Y���d:�J�pA#���~!�\\}�ڸ����K�uZ��׫RS�q��2��4�^�ߗI�0��z��|Or���t,@�1���Z��r?$�-o��ʷz���9D�آ����F�h���[F3��.�[.���u⎧�Y���U���5�����Ȉ���6��`�*�F��H��yl�*�������
Sn���.*�(�!��,Ω��#�D��A䰼@�=�@F5X�{C��l~���Ҹ��NP�ܵ�; � 7�g-����"�Qlt�sU���z��e+`����v��pa_�$���Yą����~�m|��)�����O�G�Y��Z�����+�z��2c��z�1~���9Ef�X�u!�����S��`y�Ō&j�p����3��D�Z+ޢ�@ʈ��36c�9e&߬��gM�r&N`�ܘt����e+FW��R$��N_ImFy�t����1e4߫�o/&�P\�R��,N�t([pvs�R����R�SM��[���;'��"�muc#�~ouq���i��])C�B=�$L�h��x�5RΤ����m�U(�ޝ�Xn�Tp^�y�O7�K��7�U?���C� �+Y���D�<�`��)ϮR�N|Q�B̫�w����uIZ��>��q_<<����̖
I�F.��*�I�X� O��8+�r���b���}$(�:�٠_��`u�3s��|bW�X"���<��G&t�`��5Pپ����v��1�'�_z�O���.n���~���<�7�z4)ؖ�2F�Mu����a�"���M��ǑI���g�n��($Stx��.���(��wG���:�S���'S���a���fG��▧ŽѾ��|�˿�6���|o�ɖ�����0�./���-c�&y���t0<���3��|�"�2X�x���)���v8�v䝾��B�.�JA�2
�>�∴a�y_��J��V�o,�\s�
ع���a��1���`0��ٍ�k�s���}�"�[%�4�=�0��_��>�\�@�}��W�MU�-���ڶ��}vF�ɩ�Wv>zb���1��|Z�Erv��~ѐ���2�7�Da��{:@�1�O�ߥ�7Zf�䚗7��#��B�z��w�gj%���:�&��3��*Sv�Bs5��;L#ǜr�����K8Z^�i�<$�>�EzII�]����%��6^���̨���ɦ��V5�����ò�=�o�y]�lhHЧ��ׇ�ϚE"��U�X�ƨ[��4����]��buB$��n�q
>�"H��.BS��ܕm(�'y�������R�6���k�"S�����#׭�rZ���T��yDW��S޽��C�C��3�@��s��7>�W�&��*s\`mB��Φ@�Z9�Nn�O��z�}N��T&�H�#���rt���$$�;�r=�����������_}��`��ȏ�L����#~₃�?�Q�cQ�r6Y#���`LBָ+�EO�s]�Xy��DY��jЊt(�
��[���a�_�)�7�[�j�G/����j����(hѻ��ݞ�/h�p�Ԛ���Ҫ��G�ﲦ�*�PHBe��-���.�,�����f̗�'�ݧC'�Ä�N{����C�W<�q�8l�!=��s˙�����e�opS��� P������L~�aW�=�����ժ���'m��R�@��?�ꛄ#�\�ЬxrL�pe �D��6�f�˵+��E�j�RD^�'Y�N���en�����Բ���F��k���l�X?�1zF�H�P������֖=�q��9��2��W?��[�6�-)�J��&|{;Ȍ�~���ݽ�5�p���M���ۊ�*$QN�
SKE΀Dw��<�{�a ,�'HIv��3�GŠo{��Y�Z��Hv\V�M������~5tEHh���?sƘX����5g�Կ��F�P��ޤ�%pb��&�/��S�	��v�3"��S�/H��N�ͺNf�M��'�ɝ��ώ��݋���}��w}KH��iM=;�J%
�E���Q]�.������S�#�`7��_���/�'���4`&�Ps��N�������=ހ���I#<�wc1!��d�V\ɀ�T���Kp�d+�X�J��*�vH"Z.�x��é������[�g}w�QȻ�9��$�����FK�/�ϊ0��z��y�U���;U�r9sQ���7���[_�H�e13��d���M�`�j~�;�lX�ц���
��4�"\C�9t���A+(��A+p��v�׫����n�D��,)(P��^�cS�8�kh��vv�������e�$�b��
F;�"КP�Ȑ��Lz���C%��ND�~p�Bm9�R��&b������ ���w��~P����:F��fp[�=��#�m�&u�A�9	yd��:��m%��᠏l<��c��4��[���E��~�OBCf��>�g.f�����p�Cժ'�?�S[8U� E<	}�h��ٰ������;�Z�i����8ľ�"TpI�0����!,^B��݂ľ�@�U��xX�o[���A��A�o�M!_�����N^)�^��&G�F��aM~��i/����m�s6;��u� ��E�P�(Iw���e�d��=ܧS!�!Y��[�����Q�j��&�q\��Q�Ir),�F��5�T]�B�o2��a��+gi�\+��s�*S`{$�JI��q^�b��d�ɒ��5Q,$�nJ�����!����Ҫ�_�����ԆKnbٍ@�K%����;�-ĭ��ex�.���k�!35������F3����N|;��	��A�>ǳ��9?�풻�>�O�$ JB�?�RAEE�bņB�E���|������"��������SǨի=��&��m�$%R6��`�b�%s�֭�;yk���s�D���hu`Ҭ�_��iB�(�:��ۖ$�̠�P�����ya�'�?�n�x�A���p�Tla��w�<$��ċ �Ƃ��kǛ��Mq{*��khb�eGlg������T �� .h�8 �!t#�9� 	|��&���h=߶�x�f��� ^Zp�I���v7yn�!f���k�F�I� �;2~N15��r7N�j��}@����n��!��:���;��;��OӯP;,�j�Y�>ٍ�).AG���V���nQ��V�6M{o4�q2lJRL'�-:��<¥2_~96����=W�ýJ�7��y<]j�On���	٨Z!"9@�75��*bߒ�0���M)�����l]�eKW&1d4��6�^�`j�7<sx��G����F�w�����P�w���?�&=��P�7��3�2��f�5Md��Ԅp�cr�]���N�ݧRA�o
���̟755r�Ǟ�O��<@�8e�YN�n9=����~������_��1�%�}.PZ�9�hZN��1ֈ�,б��U-�X�α�A{{�l��8
R;u�Kuf�)��'����ǡD -a=J�T���T9�8�z������}Wa�"��v���;�FUl,vc�;)�'�y�g�ꖙ���z���i�����-PR�\P<Y�Aŕ�6��%��#m�&gf+aa$�Գ���ʋ|��ܴ#4+)�ǹ�t���d�R��n4uUu�E�C!�\�9p�S��nGS�9W�50�*͗���I����P���qd����.#�}=wq�#������j�
���=��UR8��H�-����@�����(����wytK!��:�n�܋S��@A㤁���m�bL�x��u��n4)��]�6=���Z>���	�0f:�Vp)l;�;Q��ߔ�3Ӑ���w�@�!��O���qJ�MX�R�ӂ�p��ϕ�;5�<��V'�ce5i^G$��P����ܩO��,���pk8S��ҥ��[�й��	�tCF��1l[�!WS\Ce:�k��B&V�Y��)�Web�{`(A�y�m 4l��v�|��#j��z�� =�����.�5��)���v��w�x4�f��˼t];�<!P��A��S�#�9�0��ލY�z�;�S�m���:T4{o�O��-�JY��N�A6E�����6X@)*��b���<�\�=��B�y�����9�>Z0��3L�����B����&^����o�LY�`�3�P�W}σ7�}�ej�=9��~:���	Жzf�
�tE/ߐcپ�/�W�8-�?1Ⅺ��Fיީ�-��A�dd�g�8A����MeT�h�D���������OϢ���Ԏ%�G��mo����A��QO|J�Rez�\�&\�k[�ԑg���+�R�@���m��K�&���e3�d����ܜ?u��I�`�A͜Q%:����o"��$�Lfg�q;OU���upiID>-u�������1 J*{|Է@��ӻs�/�e�v���R��d4���:.N��Lz~���J0/����V	  .9 �5�̰xӇ��p`���f?��D򝷱��͆<�B��[����ʟ�9��^r�fKO|K��sPo�<�mηs����M�Au�;�7�@-MRz�k�=�}�}g3BJ^���2�(G�ۤ�%��;�`(�X�����:��,�$�'�� ��Z�WO>�Yp�O��#/DBbf�4Xl��f����߄�cP+D����x���x7�N:`r���g��DbC��/�A�a��B߻�C�q�?��Q×2�lv{
�6�_;���@a
�Զ8�X|�e����O|�c�.mzX��Z��+�c������XV+���
(�.s����࿘)�__��6M���m=����'�6��Wss����,�ngҕex(ʘ<3;����12ُ�E��G��8�WW|�P�mf�i?��	�eMޠY��/s�T�=1q���q_�����7�����V��q� �c1����P�n��EH�~Z&ux�W��qa��u��V��[0l���?qi����y�n˅A��Sj�D��0�l��ul/)sJ�+�9��9[�{®[ĪDw����%J\��J��X�HǚO�O���ǚ(^�@.<$�]�'t�Ee�kҀ�,]��L[Z�� �H���P�k��5vT���w�c12��E�Q0�W+�����T5!�M�:�k#qQ��s�L��]X��=���W;����V�\��u�a�����)�U�ԑ ���<z-��o;tq���%�,ƙ�����!$��1L #��n����HuF��q@n<��%�A��d��F�Ez���OO�	�,�Dʋ䓦J
��wy@/�_����i1m6v���xw� � �j�j�Kl����`@��z�w=���ywf ����WS�� {�oa�V>�w˔CG�� Τ�~��nK�rΚ����іB"��A<3��-mG5��t�W��֨��,�K3E��i*7����V*`z��D�b?��%��R d}X�~|s ��|=�y�=��wq/�,�߆zN���
�G_�m��	@�B
C�W�os8�������+E��$C f>����לм��=Q�狴s[^��۟�_���I����Q�!�{�s�#ؖ��u�շ���@��|�8��UX�0g�e�:)�I|*9&>�c�)"���Ï1�T*0do]���ɟ�>*0�f  �;Ju��t�D�6^!�U�v��p-�P�����qW(��x�Y�B����r8��c���f��)�V`���6/ e�.�u�3Epb6��m>r��C�3W��	�#�إ�D�1�z�������u �*����/E�;Q�|�--M�n�yMFՠ��?C�S.r]a���V��M�'�S�d�W6�Y@u%�)��;���
*�&&ϰZ�m�OUi�9މ	�v�2o#�wn���Q���-�IBDv�F� ��q-�N�ݩ��X�@� "4w =�!�fr����ճ,���T	�=I����
�xq*)�
�Y� N��X33M��"X�ԍ� ��`�JL�ɕ���$��BX2" Ԓ��|�� z���p?�P33z�)^��B� �}b�8]E�d59�)�R`	��̃eM6���D��[���>AU�V��l��.���2� ���TP�sFܬ%��*+�)?��9/�R���JEe:���s�E���NL��(��O��n�!��=y2v�0�$�#��9p�c��`���d�5o�^��.%{��ŭ<A���J�e��1���'9���}���ǳ�B�=qi��Ե�!7"����lW�1h ��Y@4�J�o�2�a\�� 3�r2u���m��܌դ3 ���}nq>gq6��6�ͮ�d�3
���!M���l�P�'�a�N�v�/S[�A�U ��S�[��:��xg��⾑.�ͬ�uُ��f��x�x�����}��n�V�Rb���pE�|1� �����3r��O��Wi(ٿ) d�T��ۤ�&��,S]F��&w�ˮ�� �|{���Z��Ilw��6����u@lĖ��G�h�$��aδ >!s�<��R6Bx_ǥ3�L��l!�w��i�qo٫�am'	�7�]zڐv`�h^몲�ek;�3�D&�=�������
 ��c}Ҡg�8�L*�NCڭ��S�~�e�LAv���×�8��3"�Q�]MSz�:T<� B���C�wu{�=�*���"�&���G2v �ddt]���-��~₮��C� ?���Zq�$����{��q-��H����R-1�u8�1�R�d��6�6:`�'ؗ+� ��]�6��oj��(��ݐrb+`�ة�&{�gf�Z�6´���_~0c@/ԅ��Gce,D	��on������Ѻ�TǤ�z����}Z]��~O�H`��B
1#g�����㥎��]�	"�]�Z����E��-&��9�&��&R�=6�D#��l�6v*��Z����������ї�ə��vt: ~��\ɴ��ql��76�\�cU�}� ���'�v�[\������W�RJ�?��?��
�B��������x���I3_죅���E��v�Z4վN�dvx�E�/%�M��N�Uw����#l��x$3�ٯ٬�s��s��P'���N���>^��%eoDk7�D9��9�M�WƤH��6o��q�'ݔS�t�u��bm�M�����X��u���t�x�tҴ�e�2Qun��q	�@�;VQ�>Ƀx7̎+��I��|����Tq�Nm��d��4-Q��:�UPa�&b���h�W>}=j�#�M����Cy�jI�_<��=�V!Q�[ʚL�9���xw����: b4X�Kf���r�cnf���}��y��-����=/�u�Ă����_�^x�I<���F(����Q�qLK\����0e>��'�c��qa����2C��W�4��y��Tݤ4�9,wV+���Gp����WH�q��mN���ƅ��L�/��!Dm �� ڋr��X�q��L	��L[�c�ь��"k�W�਍Y�������1��Q.e���CN��"��>���m�E��	�#p���d�+so;�ף�=u���x���ab�g�Ij��3v�.dT���Y�+E�n�$��a�c8c���Ղ
��'�"J�#uP8*��Wg	�l�~D[��1��O����;�F�g�e��.FÔa�;H����3����
��ISe�Gr�4vr�If;ȉ�bu�w-�B�ݐVC�=>حy�$�s �{��2h�Ki��4�k��|�i p]G�t��e���2�
`�0�9�NS�����k�fS|Ύ�`EC��~{�]�T#M�}¥C-�?K����]��A?�fJ���O��%�R�� WV���R\7G�$�-�����\�9���Q柬j��dŜ���z$m�ɑ�"M����gs�B�f�/g�N�K��G�9����i �v�江��{X�:<5��B�T�o�O��?��ExOJ�#���@"p�?QJ6�'��
ج��I6߈���R���Q��$D�2OND��U_�i��'�A:��=�t-�9(�p�[��ދ�wɼe�M��j���#-@�S�&��)�����r�xX��E�5���4tv��΅X�$��~�?ؒn��Yte(��?��,p��������Hlm(2����AAJޒ'��P�D����A]�0,��?/菿�A�� 	��Y�������
enpiq` :TI^�'8��p��{�++�"U�䂌Q]��yR���4�Sl���e9+�JvZ���~ �ֲ*�����\Ie�����yd�]b@����������!��n���V��ol֞q��a!���\f/&��هk!�p�c��٧�������pœv�^Z��7����'/��Y�U�J�O2+{@��{ �>��޶��jb>��1�Bs��"i!^�}y���S���Oc�NȆ�D3~�CA�:�Y	ؖ�1�~�^Dk��xt�K�E���s��#�U$���_�
��Q�v5ja��<����Q�F���h��X��&d?�2J�,]��JK�P�M�w���Bذٳ:�]p*�Ej���kH�����#*�?1�v�6m�<q�*/����|�C�4)dF�����s%Ŗ\��:�M�	�����_�����M^�W��)���@a�:�1աu�X� ��"���:�P���K5�v�����~dL#G��#}{���j�����v�P�|���zS?��	�2^���iu��(>��ڿ3��y]=��"PZ���`����Z:+������kH�J�	~�����,h݌�P�:���^6��Q":^�P� C�a��g4�eܻ;E��PJK}@K�+� �!����;N(�?	y�#�WY�5���ق�²��K@���� -�I�(����7�|����ؗA�-���Eʅml!�r���?�5{���jh��P~� �� ����o&�,�t�kS����(��L�X�eJH���i%�xF6��x7�M'�LK>VՑN�M�(ٰY~�GaӶ��hhz�MJ5���ah���.������9̕]v
P�y�,���@��P�c6��)T���v��6��H�*���|�M��]���W��4�gQ+%lK�RaK;������B��`�,��ZXZO~B��kK��i�o�p��1y�g܆��̔�x3�a*��I�VW�j��}U6D�+��/�S���@BDJDd�2M
����qth�6?Y#cϹ�ut��C�Ƴ�Q��fF~maK�Q�>�&T�ԣ������L�2Q������� +t*�"(?v&���Ƀ�G�m�D�4o��!|8�|o����A��wv=F�aO��?p��ԅ��E�}�������b�}���+RVA[�ꫜ�uR�����{�B�"jL�(6� A�g����/�`�w�&�'� ��Õ��
���˨C;���FMΥӨ���=AR�A�i�`����X�^����g��s'�M�7�4V*x<P� �KtZ+x(�r�JDܿ0����ji5�]�8C(�A��%f�-R�l�s������1�o�!W ��{򬫱l���۶�^�W���hr	j.��U9�?��:A��p	����[Q��!���3�)ɟCD�Hب(óA�^Q�'@P���l��fTV�
gGy���p�5*Y����
Px�i&��ҹ�� k�Sm��p��m��������S�غR�/˩�{H�"����riM��ϟ��;��Jo����?t�kIN�~�+!O��\:)@�|(���u��,�쎠�Pc}���v���(
�4FP�",��xz٪c!�oϺ�n�h�hT�(C潶��C��Ȓ���]�x����5Ǳ��I�z@a�.͆�ɪ ������Լ�g~�nY��ERe���]j�X;ڥ�۳��W�GL�4O#eQ�:q�nA�@.��`f��g�q��"�ګ��3O�~�z�T �+#
� �mh��$�ZJ����NXE�E;Z|�,����������V9�=�~��,R8e��Iu��!%+>�s_�UM�0s����epo���cpA��xY?O-g���v����WG��g&|�k��f���5X,c(4
�|�s�ax%R��L�/o���1%o5�A�@�;���u5&h�t����)����f�"�l.�)��b�຤��I���].
ٳ���{� ���]�߻b�4Ug�ި�)45�Ͼyt8Q�A_0;�G��|h��E�B2[��O���m$5
w8������r��ˋ�~0�(S�>��Di	�]+���A�� kk����u ��h����b�6���	m�Wp�n�-�S���_�Ƌ�����d�ҁV5&-K�c�A��DMx[���}�X�c��s �/;�e./=�oWeV[��r$��˲���i�r����m{����֩�	�� ~�Mr�H�ƭ�ݴ���{�ع�f��K��$���5a뵋��%�_�wO��(rBB��Nu�Mb��z�a�VV'����5h���tV��@����n��Pe�7TƯ���RbK��#��_(�{�[GM�p���)�t;�����=��j��U�z�9��9��3��m*Ÿ�{)#i-������ƽU������؃����p�*;w�)��1s�OA�;����w[!6cN*E�`[���ޜ��M�y���<�'��*3Se��<\㖡a�d/O�������@t~#x�u�edgz��` ���8C��<�+&�y��X�'>By����ψ)t_4ڏ4q�6�D�a�ڗg��?vnV����3��G���&ܶ��V��?*�2�B�Ȃ�zȢ�7`��z���L����w)��h�m-y=�4�������۹d���4?� ��)K��V����u+Y��Y)��`Įޚ�[¤:h��t��~����G�I����&��"W���p��$�(�È�j�v0n9����6Z�S���'�M��}V�~�=pt��b@��|��Fg�mc����,����W�
m ��A�"U��Tj��,hT]�nT.#w�I����=Ş6,cI;<�YOHK0�W�B}�8�%�t�Ԫ�o�B�����q~6�zvpjE��������WO0j3�$�� �-��4"	�P�4�%T�[���NV�_�������i�`.C�˩��j��Գˊ�?�Վ?S�9�3����H}�v����	��q�$آ'�vQ�H�.�J�a�p>2x����FI�������ls�o���p_i�_Dyֱ
.ꏍ�����&�{�{u�A90�[̀:�;��5�3Z�Z�L���W�N	���3`�r�Ի5~�	�>���� !)�- m�/�z��B(�m�ta�'��S���O�Ȥ6�X��ob	s;��g<�(�4Rto&|�����Kx3�e�	�[]��K��j	��X9�o>��]�����&���u�,1��3s�����[�$�VCa��3����
�#DiVY3��D}��0-�&��M.m��v!~���S��$��%"
'�Hg�D�ݤj�7vN-
Uc@��y��]��A�S��=��O3�����폍���,��T��9�߷��rIFlY��w� ����pf+�iPm̑Q� �,;#�q����E�6���M�k�}U�W�ax�M������������n�&����{����m�e|���?@W'��
�t;�;G�V�hKƛ}�W�d�)�	�0^Ƭ$��ʸ���#�+�8F<�\�ߙ�w��i��6�#�e7���E:�����}n� [i��c��P��;��QY~��r�V���l�7�q�6�������Vc��������5���m�� �k+׎ʉ�MQa����v����L�{�S6�_5��8�¯(�O+MW��Rb�M1:;mj9��/�sF��o��n沆��̦>�tw>2���~6;�������0,"���1J4�嘇f�_�����,������-c�����
�RO��{��ן9���ʖH�4��N�nS�xhc�a�^2D��g���2Q��F���J�A��0@�\ˤzL$���WY��cV@|���Q�WO��=+TZ[7����#\�l�P�w������~��G����c�y8NΡ���(yO�4�S��;��1�_\׷%2/�=���1�Pc��LUB��w�/T��(o�=(��SM	 ��I*!���|木���]����2��3�7y̓1��'�����������s���ۢ`�ٯ�����Ms���'��ߟuե"1��{ A����]�|!o�@�zX�jl.6$M�C�����$1l�.%�w��p�p�+�:o@��V^��^�5�%��~<�ch�����kDn:��Vb�LR�,�+^�)��]'N�h ��J{���f�l|� 8lH%籼��J��U�L�m-��0z�p��d��f9B,��b(4�wr�۔���&�z5}��o-d��89�!��P��)��yz��`M�~��R�� ��(#��>�D�z}� j[%���ŧ��N^�t��X5�=�a.L�C�E����qQ�_j�)"N��o������L"��`���<,vQO�%g�����m�&��`�Y�A����CF\�+l�"�X���(3�=�t,�6�v��mB��?�d-�`��RӸ�M�+��Uak��S	�+&�~�3L�z7�'䣀7�M�30`D`����7CIe�\�|/�H����Y�mK����s`��Z�`��p�u�g2���2%�i�a1K�	Z�����n~�h�S�U�&��y�ᚌ t�#�h��j��s�c�ī�P�@S~�Z�t�!v���?pN4U�y���^�������}����3��?��&����Zm�tל]�A��X�+Y��L�y4$�dX<I��_����l��R�nF��'��������m�k��|�E:d>�H]0
s���F��]:b�Y���1�"QF�nrc9��Zߟ��˷��xW����Ds ��Zg��_(q7/x�.ߘO�k&n"�?C5����A��L��:*Z<V%���Y��V�c�93��!Q�d���{��q="K_F);�*Kc��3�HC�Kx�b��!�b�.�+D����$��Ϟ�Q��V�⺿)?�3�l��A�c�8��w����$�{��Z5"q��d��aî�^W}�բ����LE��(�w��JJd�8=�4��,�y�҆A�X]OɎ����;�/�#A�I#ڒ�t7���n��C�v�j����%m{�,q	��b���a?�#���~%�D����u�������b��y�����I�({F�{��kiA����&M�0�/x��7T��X�i�\v��gq����m�|��^i"K�GQ�<�9#��i��g�q̟,'�J/%�ٍ�$)��W��uvp}��u�⨼�(����ȿ��w��6�O�q��jI9�и�����.m��<2������^�[�Z�4����9�?���*,����B��JKLV\r�Uc����*�|��y/tؼt��A�x�Gy��ڬ��,�T[XbEM��U|ٍ(T�TW~;�tSD�"%^�𠄘�Uyp��Z8c��`�� UQ������L�~��ɌK��/o�A+l׃�\1���$��mzjK*F"BL��9�IBNDVݿ#��;�F���f�u��YU�]����u�RM���߷K���M���2�Ζ�.6�w�@1��P51_6V�@�Kt�����cZm�u����>y(��굏O��f%gUr/V�a�P��W�r�Ja��2�%�l�$z6���\�a���f��\��E�1ƕ=s�`s�>�R�ނ��a����$Ϸ�4X./�7�8X�?:?��-���,D?׶����3x	?b?	�n�"��ǽ����ٲw#�j��+�8.���O��Ё��Xn/���h,�\�s$5<�w� �P��]F��1]��O�����,���	?+�g=����@]�����'�}�a§:�y>O-�e乨�t�T���J�Y�h�Jk�
宔�E�P�q�~Jh�]�d5���E����c�Q���&���X�����gD�R��f����~>��,�-�o�j"���`PH��j!��#q��I���B��|"a8�'��s�m�������j�\@-��\�=�@:C\�Sr�y��0E�@Y��5����S��-�
bǦ�����l�T��`��nMZ��\���N�&�DjI�6n�'A���~Y"at���4�6`�]���s��1ʢ�hU�x�Zp9��8�T卑|��|���G
���e[��G�N���^�I61N�$����lՏ@Qj�V�^~���Й���K���NWG��$�|��R�#,�����w�Y�x ����c�"�P�'%�Yz.h���}�s��3�^6uP�^-;Y#Ϋ�i�C�쎍]���fd�m��n���7�v3�/f�������닜�Z�I���#�;��k����D�	�yuӤ/��!'�0APojU���u��?�^B���R��'>���vA��E�H�(BM����7b����ݾ��[�Ȱ܄��8t����{���a�KqEI�2B���C;���C� _[��������`=Ev+Fii���uYE����n1ōd�B9!uI< ��|-�q�[3�D[�3:"�i7�6�8��^̓qc7ɯ?�jr2�>��D,8�a�vU1x*� ��qK�/e𾝮|aDm�T����H]8�+�T�����&,�׍q~��?l�W�H�~�84��T��Yh�
�3���&4�ț�M���}���{�j�S�8�DK�LD$����#�y��| F0^��TYt��7@�~�x��CU��݈�՝�ĸ���33p)x4��b�[�l�`�#]���Eb&�O������t�%^����Q���COP�1�����M�� �`*�HM����t:q����O���A!u$;_���� U�k�I���$�XJ��_!� ^�e����/�x�W㠃�<�Ώ[�Þ�.z�:���\�׆�lKtz�<���kEe���Gѐ+ ���M��L$k^���)��e����I�<u<K���q�P��]�y��U���7���h�E4�{��ay�s�F>3Y������< 8;ՙ�gێ~BO��c" �ђ:6u?�z{\Z��IK�I��f�U��.\��O��Ooݮ1!Vsm�`m@��a�e���7�>Ο F�ló9E�rf_����f�Q3X�S���M*���{LX�c*MyV����B(U0��E*Wnr��76�1_��	�eҳ{4�L��p>k��eԊ�0�-b���08�Ԡe�K�$�*C�-(�L�l��.��,�1�TOm1��{R,��<V�f����}�XD?~w��L�ZT�q1����/j��ǉ$������'tOaH��	 p�zg��R��Xm,^C x�������(�r�Ѧ֔�i�o
�d �]��]0��9]��}`6�7��C��b��!��
$�+q�Ya��֔j�u,~{�|RGh#J6*�q�$Rq=�r3�TN����*�5UDyf�ʺ�q�:i0G�(�NZ��4n~�CfO�q�㝈&�5��s9(08@{�C.�/T��3�P��!�][���m��7�H,�}P&_�ƒM���Z"`����p�0����`��m�]�}_��>7�q�V�!�)��ώЅ�>亾���ᛊ7�&8:�6��.��l�ǲ6ۼ�	 C�{P_�<��i��5�r-��Ӗ4y��>d����K�e5h��'���k~�1ĊXg��/�/��V���$|$/:�1��I_��:�s��^U@-4Ac"_\�poW�S�],�g�OuO����jѓގ�AD!����Μ5w����U���<�䏋�����Nb�!�|�@���D��y�����t���(/��fF�WWi,�D�T3��C��o`�~�z���R�3��_�]�)0��nҫ.��3���$��7�zHgS�oGxRJn���]R��|.;��dh�q�=�,a�J�i�>>�1�
�p�׻��=���Sׂ׬b��T@�y�Qf��|,��q�+�^۞L�k�Q�$r���
0p|y�ď8e8��*	v1��.�˧�&ד�a�ĕh��'C�x(=hMV�g��7Af�N��ɵv����w4SozՋr�{^�w�o8�� ��oq�x �k-|OJA>��7y�'�Jٞ�����U�+��s[T݅��[��j+�@EK��:���_I�F��D�ŋRn��ɘ܌ھ��"H?��/�ڽ�,^<B���KFZ�w���̉]�Z����կy���[V�%p<O���8�Ȯ��|�K���F��l�=���<`(�E��m~������5�`�b,?J86\�4$��H=Ga��!�H���=6Է�>&��#�a�I^F�P$�#@O�D:��:���q�8�.�6cX��R�R�2?����F�"��@�� C+ϛ�n�=:��v��z���q�Fa,w��U$%2X4�i��x�������¡Ce>��m7#���s��@������t`���C�P6yb9]������9�f`�e�5���<(�Q�Zb
���0�M�����%�-M�rN�z���'�BCv�-͇[L�S��=����Y�ˈ�|.E&�������#�a��D#Hk|{����.�)��9�xj��G� p��!4�&��T���Ӂ����J#a�t��Io�9ϡ�f��GW����g����	�"N��'�$��H��}<���>�G\�Hq���<�V��Ax���-mjt9���v��&�
HN<�Z�KФ��K�hT�V����G�[���N/[ںA�9�|(�Ƈ�T~��ۥ���w{�~���'�;��͵[f���Rs������cL{,��(�,�'�W2�gӐ��:G8��v�G#h�����n�hR���[�F.X�P"��@��p�<�uk�y��OEFBy_9W�n�V�䏣"���J����oS\i��L�X�9x�����=ϋ�ޝaX� �����	l�_�.���A`��!%���g+S�p^�k�$VDs]��A9��5�4���̯@M^N�.)�9���޶�ҏ�(	L#�gI��)�&�in�n�\  ���V�P�������]�5�.W�s:��l�yا
�幷� �j���ѵ����.�*����&Rs��r~1x;`~6���f�$l�yۍ��;���y	�[g���$����#0tk�����	�T��'&��M�2�َ���{����<�:G̛AHY	����'*�ᥞ|�)�Eٓ\y�.�O�E]�?�.Nt�R�<����5PT�OD��I�8<�3�P��Ț�����)
����\<F��K0�=yv�:��-j�n�dr1�H�I]q��i��-���\Ӊ�F��H��*���x���߱��� V�(���f[0�j��,E�o˖�FFp��t�y��U)J�nz<u����氀���e[٧�)w�ډ�S�KЮ�L�<p�K�g��ʆ���C��l�$�t�	�掮`�4!��Q���2����톑�Q�&�&����K4Q_�%�.��0��mG<X���}^�Mb��8�|�^D<�l]#����7k�}�_AWx��L�}D���@��_4*'nr������0"��d\�Ef[8f�?>l���N=I����.s�zS����TB��D�����D����qX�uɤ���@���Yf��{s�[@� �n�`�إ�b��9�@Z]꼔��H���{���'�h����o�\���Һ��J�|E�o�TiY�Bcg� �uS��ڙ2��e��3�JO�Z~ZE�u�NA,Z����b3V�5�� ��92�2Jf���)�;5({)�؟�rf�g�(x:�6(���<���	,�N϶���b����d�;��w�$#��Jp��9z3����Im�D�r���7!����N��+M��g�L/FU�����4 �>��tA��J̱A�ʣ �s�m8\�-0���pPB%A�m뢲�;�PC�b��]` ��X�W'��H����妦�L������9�mDl��Wz�z���NH��evi������\\�Y�F�����SK�RΉ�ɐ񔶥�^��M����ߘʥ�{}OR_mQ슛�'��|�+�O�R���Ř�jJ	.A���u�k�h��9�.ը��{�s`�����aàp)R�u�}�m�í)#t��bΫ3>}�<-#���x�z+�a�
m8O>$ ڂz��c�
H*>��������`��4���9��5������<	u�]��(0�W�Y�F!��#-_�EI�O"�gKR}/lv��,�AC)9VZ����
V���*u�i�8#'pr"x����|���$�c�<o���"�K'W(,A��Xr��|<x����= Q�{}h�ǜU�9������ֽps���� �z}�ŧ2�rF �J0���i�"/���(��B�����������'4+7���@K��jxG]c݁j��]c��X����A�c�1�5y����s�m���#�.l��2�J[���s�j�����&t;�۝h��.���'��W�� �k�l��$�b-:���Z�v5�0�l�@������cS���!���[��Ğ5����n1cN{��f�F���z%#��R`�.�kR��h���\����F��i|x����<����NB��l��}iX��	�9�N�K	�`�='��-9OE_JG�k�&���%<d�ѐ�Cc�����T؜H��A|�#�}0�P;�9�/�1�t�u�)u����upq�������{ ̼��Y����DBPE�h��heؑŇ�޶c%�}L�d52���}�C`�yQ��x-0�o��cu�o��+ Y�a��'�x��,a���5�P�f���tNO�q�����3m{<��15�{&#D�sg��8���M,��]u�\���9��w��NQ�1ɶ�mQ���O�pa��~m��j��f�K�^����B��ϐj����p�G�9��iQ! ���6��>5�`�ҝYhNt���GE���/��s��%	�/T2_Vjug,o����xuQ�7�����s[$_y�ڜe{"ŋz�s'����fÙ?k"ˀ���N�[s��*H�j��&�h������Vʞ�J�/���_���ݐ� �O���
0^�/@k���e�M���0���ef)@A@<S���eo����Ah�+͌���t*�ԲTil^��k��+B��n25߾N���1���Ǩh ����"�8V֣籮�3���ꃑ��aK@ǆ�>�#���kz.;���`(2�"�S{
}�ɼ����^��!)
1t�v^໶��h�f��K�a�,_f4p��f�y�,%0��/ɋ�_�K	�P�]�"��i3	Xz��Z`ذY�B�K�>��D(�lP�'ɨT�J�&�L���{�ԬH�n|B/�g�,��I�ݟ��Ň�W�������؎P��ާ	0�jeq���꯵+E)���33o�*^��yM9��d��t�#=[�#��x*��b�uUG��j�j1�9r�)Hr7�\�r}�z�����}П�*?;�@��v����-�����L�7h-a`7���k�_� }l��⹘)9�<i��>�m҄�Z����߃�ؼܺb"�r�e#�6?�]� &s#��C�I떣���u}	$B��Q�Q���[,R[{�u�9e
'���h�[ሗ����/-Td�#�����h�!�x*fvH3���^Gsaʳ�%|�`�Sr���D�D|�+��o��U��V�H��6�����^D����%�9oi�7���r1�pP�/��Z6��'�]'1������Y@r�����шɲg=R�6,o#x�/1�㰳�����a&���"���+3��E@5�_B��#<��}��=���<e<=ǎG����
��	E�5�^��,�X��������I��Q<�<l���>��P)ȧm"y�V9jK��(:��1�>�*��]#����G��(S���m(�Z�~�ө��gf���'ǧ��@�?o���]Z5V��L�����p9�Gm�g<�`��v�.	�i?�W�Y���KX���#L�lZ!NZ���[��2��yh]��CgQDu����p=�*��&���e/�T�d�p��B�#�9�:p�ڶ�Y���lӥY�J�H�����X>(�VV�T��r��>Բwm���	�s���L��A�{-+߉65�>DFRd �P5CLSH%$��gD��L����D��)����s�é��3���<!�ض�2���2n����W.�|����[�0O8����D�����8(��j��n��H�b�5��W�Ҋ�����
�Ԧj�c���:��������h�
�E)l+E6y���2U6M�(,��	�>��b]�Eԣ������cu�(�&{y���В "i��
`�\���*����A�o>�#��Ԯ}�C�}����L�
�:O��V-� h��t�c��R�H�ez�%鏓� W�=��og9�����G��1����?a�Ul��ݬ!`4�t��>9��7<�`C�D�_�� s�,=ې����&Wi�k�#�Dgϳ�n�gu�.��c��yZ8��Ox��T�>���Ğ�|�
��@�T�Jm7C��rR~Ҏ��s�Ψ֎jy@�u�b>,持z}ѐH5�>벨�����v�*n��#��Ҵ��x��gi;��x�V��҇�7,��@��󫬏�f�Ɲ�=��Ł�W�+��18l��q���l������z�ƌ�))�g+O#5Pg-�n�_x�i��������݅wY���,���Mቀ���q2TTx����<�l#�*���
�)E�~#�3������G��ӻR�a�ۏ]cݹ$;n�k�4�MXr��``ߺяQ��=W�x��Ok�M7y.T��>%�Y׷���0���^,��7�H�i��|��[��Ҁ��.����<d��=��\c�����E��(��+��)���=3ó���DL�g���D%�eC�۬��z�4@-��mU����2�8�\ߦQ�Ɣz�C�e� �a@ۙw�udOwcy���m8�~��3�tRHSp���[�M�B'���O�X�� �@xM�h
̍�{|TLI�%�{Ο�r���Ff�4�9����F�*�[p����*�����O��}Ъك���,����튊q�	7�����+ g�*�Մ�E���]�)�Eͱ�!mYؕ�O���
���x/�'�^㠚К((��g"\/�pJY ��w�2�-�s(��2&V������~�ԛ�F5E.����ż`�W���!%$��b4�٭팜���ۘ�_HqF��t�F�7S��U�������&x7*�o�>Ql�����H���
(��6W�ƃk�
h�g�j� ���2'�:��x�8����G\%��g�&��s�X�s�1����W>�jR�0��0�']���X�!�*����"C�J)�]��p��3g����0�q���h�j�X�Yуt�E�fs>�k�J���M��Ҙ<}3IA z���+w�t�Lճ�IH�^��_�����J���~[q$�ȷߊD���T���N���ol�<�
������t�7�H^�<���Jb�ӄΓ�{���{��rlv�G�|�h��_6�K^a��)&����`��!�h�#�*-9�����g�X�S��Τ�Vv�sS�+T��D�YIo���&���`�^�����.VY=6*�7H ߸:�����v��+�����\�^�,����$�s�b�䦹���x$/�.:~�E4n�K�'&Z�>�P1�\ό����_���gDG���64
 X��^d����B<�W����4x#D���yC[_YK���RR#�^�m��&W�s�F~�9_*�Y*������%oxf�P���f�B���ry<�]�n|U��E��If�@�����b�k,�e'ROVhw�ٻ:����0�ABIվ�P��<;���3�I�&��礰�h&(�QU��5F�2:�T��4��E抋_zs��^��m��r�*�a��_�A"CfN��n������M�D��a9�+V�x�Xj_$��Giov��Q�f?�[�.|z�U%@wOF�d̍e��4�#㲨����B��WY<��áv�LP\��!ޖH� }7E�D�QS|�
���{zHw�}���DV�r�e�)�#�G�D`��۠W~��Ǚ������^sf*.��X�pr���Z�q>��A3`�~��U`UMP�j���ߜ(ޣ�ɿwD8��B�S��kq�� ��I0�l��;[f��P@-��%��:0�JYq��=������4�}��Ul3x�R]��au -������@D���汰��J,�}����eS^%�2��O������1r�f����K�Ǖb�L����7s�!v ��ib�#*�ę�.La�G��.�X:b��va���ا�-�t��7
SV�廝;O=+�D>B�7[R�d�ח5��U�Yb�R�a�\�(%ݙ�^7�]ո&�5G�'&S�&E��jr���6Z�)��1�|�bR�E5��1�y�R�j�k�}��o�̄�"1  ���f�u��uv&']g��#o�+!����?,��s�k�_؝qq�����UPIA���S;��uwh����'4��AY�}�[��p�w������)�R�(>1��v�Vx`V�mڤI�arۮ��>��K���IJ���o�O\vU$ry��	�}�!�J��GF~�."
h��1�Ze!V�������R4��Jɦ��q�䳌����b��^aɲ>̌&s*t�w-*�L�>ͫ�g�&�Fx^��G�f@`7�`�C4�|����B�u�Q�:jy&�v�9��rd.懒���@�a��&e^-��(����  �m��	%���7'0�q8���k27;O�O��]�W������-F��l&���S�� ��֦�22��X��Uh���D	!��KX�fxD.��{ޒ<ɻ�=W1eN2�;BD�lU���C XN'/����²�2���e�=�Ueu2���F�mNm�T�$��$�\ޟ��<"�wYS�N4:��ff�;���|x��|k㖭C�d�z8{�i���
�O{�n�X䯢�5�
�\��w��`���@���
���2O!g�iE�b��f�W�W�ei��K������H�g4�h������v@{G��E`�	.����a;���H���b�;�����KjMd<Oغ���X!�ާ�7_���gH�o����&��M�_����`�� [S �&Lz"s�{ヾQ�bño�-�!�2́�O�!�~���~�Y���Q#�B�&7��Ҵ?^@���)��Kw��/"�r/�#؞��)����@�釪
{[�>�	()oJ�濫^�z��;:����-L��GV��U)�|�ޤ8��
��6��f#��	�1
�S��9�����[(GC�Xt/��ro�O˚X*^����k��76�%3�p�ˁ/ۮC��j�a���#�o� [�f�bZ
�Z�
*>
�2 <LIr�Gr�8x<ju�!<ZX����w勳����S���>�J7x�&�p���12OOp��|�@��m��w<[C�ƅC��Ψ�"����i։��+Gu�\o�] �j����P���M�O�(8�������F���+��m��S�ro,�k�vY������;�L$$�h��}\� %�=��Rs$�D���q�X��X��1�+81C���k�P�#�I�}p{��1B�.?Mu�^ͮ�04�{6l��Fi0��\�=^Z�q"�z��h�����z�v�1<}�	]s��m|�ớ7P�4�8�:�|�fG�R�_�$��t�m�����D��ٜ��ЛS��~���L��_�E���_�RJI9B�7����_�M��G�6�`{@���.D���h���Yʋ���gf�~'��T>�qaLz��e�)���cR���ny��0�{�ݮ.S'��QQ�w��}�q����;��L\@q���m<�x��iս؛`�?�3;NH�sH�辶~��V�D�E��ѽ��y]wa\��ئ)��r[]?E�+�D+��;8�l�F�y�_ߣ����u��h�\�xngo��-��]K�p�n�����~Z5:E}0��I�.����u�ھ���VlS R�<����*e�_�8й��wcxQC�*:����Ͼ'u�O�.-'\Q��%0N(�z	�����*[b¢}.���,� ~�h�<�ݘ�1`.�)d*M��@�<Kc��{��V��'_��hG�r�I�H�t#04P�l4�ѝm D�� �:^)'w�)L����c9߳���!RE�<�p/��c��X	�h~�:��-���azV���#��;�x 󥮦�.5u���M^=����+��o���>2r.�8#�S�Guo���l�Gsw ���wZ��T�⏡N��_�H����VOff�
�P�1�_�pFz��	(��,4H3�qҚ�\*�BA~��q
$IZ����2��X��vtx�O�Va�>E!Mo�P%*�Ҷ���D�'�y�2Q���vy�	7��T.S]v��_�g5�խ�<�D�l�6x'��*,ס;�2�ܛ$hh,�ҥ��@v,���������:j}�a�#y�Z�|P�؎�!�H���p-~c^p���馷G�˃�]�0:9,�6(̎�Dv���{��?ٞ�@��a�B���ؘ��F�ϩN�%ܧ�_�����c�3>��D\���|,Їm�r���pC�G��~��櫄̱��DD�� �E�pt ���C�^�'n(VW1�&1�U���0�����\�f�V��9�k��z�z����ɴEW�c:���y���pL�ץ�k{�=�W�FpJ_'[a�Ah7�;*.^��,�,��w�_��7
�>���YA.j�	y�p�O+��"�>Yqfv*�3{��C?�U�q!�����8u�X��}Ռ�*V`SWL�Yt��559�ל&���V��������J4��o�V)�:�~ߗ��w�kF�-u��j�qh>)F�sdB�E�߬�բG�Ƭ,S1)-���oG��:��pM*Ҭ�����l~������z�``�pK%w�p�R*�<.����|���${0��)qi��z&�{G�Z')|c���O
l����|Ǝrؗ�jg�J"�,���ǿ5&�`�1g�&����#�^��� G�>%h�0�����E�z��8{���-���N �m�H4���W��Ot�A�������E�U7�SjW(���[�����@o T�2_WU�G!��ң�����U���(�O�Z֪Z��"[@=]q��[C#��4���z�͵�=M'a��;��`���!���ЛC�x�KFYY1���Lǩ�'ׂ�Է�^|���u���*�|�[ T�Z.���;��@mP�z4C� ,�b��gg����x����7����x
���aY`�G(��3�5Aφ�/��Ű�S���ܻ��9{h� �eB1�/�3�>ǃW�-m��ґT6����!��"E���=A���Lb��i����l<{��_���QM�������R��{N���D��
�PJ��ZQ-�L��Q�-:Q:��\!$�Nʶ�4�7�S��[� �Dl!��uT�7]�k����Y�g|��4澘�m��s������jp�>`��y��Bx܀Xij�>x�����.��#���3U�`��tx|oZk��[���yz�iwd�#z�ckj	��$3s��$�+8�{�sD~-9J�4�o묎�?�͡`��I�6h^/���ϦW��"J�[�2��]��-�g�شm�$m�5����;6^�hiu�U�Lb�U0�NP���e�$삋�W�>v"Y��y��)��Xh	�����
Yĸ?�2�q�n��$����٤`��|�M	{�%����z틗k
����N}pB	GJ3�"|�[�}�-v"~%���p{�E���W5�5���Tŭv&��5��"�Eb�Q���t�VA����P�Ƃ@���չ��Z��e��D=�Id�$��!����k�ۢK�`�{]�l���Dlz>.��2PB,{���(��7}ml8^�N9�P���3UZ0j��
g��(�o�*�H����?�����e�R�S"�G�%�2 o�4a�W��"U��Cġh/ɠ��D좶�w���uvW�� @��h�m¨T�+�TmP�Y��7�?
'Z&����A���(łev~�J�z.y6wz�I�[�6'���V�"̵UD�ګ���� -i|{2�eE�|��x�6��R*��X�E��޲,WrgER�G3�Ϧ�^������� 
�n��n9�Q�+�r��!�A�e��R;3����(9v	��!+�z[*����/Wʰ�fT���^��pQF���vv��fV���>���3��z�\�8��$�ޫ�i#�4�G����A������-m��q#�����>#D�s���R�k(Q�/5��nFP*lt#(��z�z#�b�.��H�.o��]U�0�m�%h�d�R���ܫ�_FX@$nZ53N��P����-�oC��_Ϛڰ?9��:��&/��oo�w�C�0&�w.q��尢XP@,��E
�BҶ�(�^^B~���g@|U�������Q%�;�Ι� :YI��LI��%�=s��`}D��VA�'�� Y�~���Im�-�Y�:^(�rts�4�~��7�@Ϋײ҇��\�R�95pem�Ht?v�(PT���&9�c6��pj�-UiO�KX�_ۇ��0t���X�8~���������D�o�������#tg�w9v�szt;lyPК&(c��m+�U�Ob�=���u�am܋�kl�'�\�+7t�2��^���W_Q���ARL�2jQo钷����]�����vǫ[ �T��0<��x�I݆���D�uB���ҭ{��r�-/�"������_���=z)y��;d�W����[����w��p�wL�chOIe�nzL����d��=��Yz��?|�َ����{��~ǃ�2��StrF���D��"�L��qg�=l+��Ti���>C�ao����p��Dд]�C>�X4������"���e�B�o��T밆z1dң@Q����fEȕ����2.�-7�א����B����D�̞vb�$�䃣5Ѩ�bU����}�?D|�
����H���bf��9������P�����>()���C�Y4>D��}7&ï����r�J�N;�U�g��%��r?ֻia�d��b�α�)1�.�h`Wf%�������-#+����q�-�Ax�{��CH��H��(���
�j'oc�/��]O~3�4�E�$�ސ���w"s�2�ܝ��I�bZ�������RE ����p�(�Eb������g��y�I����d���5�v��5=~ww�a�CP��8#;6�U,?{�.Z�Չaך'�,,��Oor�O�-?t0��/�4^h-hC0&�*L�intK�^��.�m�����f.vz��aЊ5y�낑UN���9�+ı�e���N�	���P��{Y2^�|�4l��o]E��4�T�q���>�[M����{��%S�	St�8��ѣ�]J�
�E��E�喼.qo
v����}�`B��ïn2"B��&1�Ȧ~���,�>I���qWۄF�p�8�/��i/|� n.��V�
��B�H���h(�OD,>�:F�X�v׿Rn-�Fp�C{���a�6̉�{o��X�{۟�B�@���#��*I��;4� .��!ϓ�!iF���~5�aO�u!��yf[W���%$' ���M���oj�G�葷;�B��Z<�a��k�׀0�����
����4FwvT�$D�[����R�4X9(�Ι�@_ `YR_2L��=�
N�.C�"������/��nZ	��꣫�f�V����=(�V17��;U��l;:�m=<ߪ�	�(T�E��	8�$|C��B���z� ��ۢʴ�Uى��'��x�a�Z9�^òl�	�8��č�Y@_:��8�Y�/�@�����:��+x��Y�����,p\��T�%��g��J66׊��S�C��˒�Ia��n�B�3΋'�=�j*���6
h�E*�VZHo��z��2�
0Z ����X�>RWq[T� �)G�O�`������W�!�0�Z4Ax�}�3<�# R�����3�#͂fd�p�^4�c��-М'�K^v	p4�	��K��F����O_s��Ep���䈼'�nX�<��ΐ@��6��Q��1���*��q���RO]elL|���4�2��#[d�>��~F����)L�h���zf��@�x�<�9ܱ�
y�a�wa����Y�}\K��J(z�!��zUv����&b�����n�}謝'���؆�$�|:�K){��I�r�~�I 7z/���L��\�V_��	�Bak&���o4�)�C�|���N��K�oSe�\�`�<��%���ѯMI����a2E����Gb1 �������	5#h�x_�Bi��Ȉ7FY�F� o��ϫ $�c����K�-MW]��⾒�s��n!TS�$��+˺�8�gh�?�|M��j?��qp�F$WS��	d����m��+"p��ֽ���H�0��$���pFOdN"~�-7��r��+������`ŗ#�@��f�n�ҋ���c��W��\ֈ!�e���!k0H^��M�{t�ka���+�}
<]�_%����{0 ."Z{��sL�0�T�}|��T�<4����nD	��֕U�R_�f�\�l�f5(�E�Ќ���ٽ!~�=]�bU]�}Y�܊��M�[�tix:����|/��g�X��W�_@]ӝ�%�sJ�u#��8ę��M�
S ��\����#�ߖ���(���E2�y��ǿPנ&M��������H�^�9 8E��.X�Jf�+�$���0ӷ���c�)������T�'���ڣ-�X�p��#@�v�o�;�~��GL��.l��%��\$#�n��{�W��)[�o�<xK���+2ī_q���Pӯ�maV�w>��2ט��B���t�7+{�Dwn�­���|ؓ뷼�a���8�an��n�i�G̻�|���)fyz�Bn��m��ˑ���ȣ�� 1�w݂���7;$�O��\!oKأ�؎��o��$��`[p=w��C��N�I�)�dx���MN-��U�E�<W��3�_��W
ɛ��@wZV[����y�']�|�i�:�DD�?{�}u��޵MIJ@�����@���A��ċz���IU��N���pF��F�4 �4 ���8�t�$p���c�-�N�5� ��ٗ{�Lk��m)��r#��[���Z#�<xu~k���gq�Q�
�r���}z=-Z�ٜ�g2�3U��M��|c�	�'���+6�[IpQ1�@�cE�:W.H-r�UBL�������$�'"��o�\\/W�
&,����ʝ��0����^]��� j9Yܚ��=��ѽ�y�4�x�0-,m2f������,�� �Q��񎡡�k5�j!�Ȋ�n�6^�S�]r!���%���uJփ)*C\w^Q��A��a��b!�?F4�|�u���=az����am�>W}�01F��J髮��xg��U.�`�Z O�Ar�˼K�[�8j�0�($��_��#���c�_ތ�~�[3-�ҒU����CcH�\���*�k���JjF�CK&+Bܨ]n���G�g������Տ�4Ĉ��h�<�bS��!�n�; � ��y���c�`J�gf;���F�u�B���crJ�x������ԫkx�4�1Xt�W��kF�O�s���)�0�>g�ʰ�����1� �^�a��m�k��h�vx�ӳ�p����@@É]�8~L O���� ��V��B1;85�_�{����{�j<z�Z���},u b�3��c�.�\d�59�${C��S�w�/�Z�=���@�$��=�V�6���(Vz�]��ϩ�k�������b<��!�"����CFU���ء�jd)������X����l@�Y��v���|�a��]���	/Kgm:��a*�3Efv�žs�2�`�(�~|5���2�g-._�f�5d�2 �:������DI�;ٍ9G*���_i�$�M4�!さ�ՙ�pP�T>�n�X�s��ȱ�;��{E]ٸ�lN�r.�ˏ��℔��Ȯ���/�b��T�,Xs�s�Z$k��MqyQ�]�kj�ҡk$�K�.���{��;��>��b�QUf��?.)0
Ħ_��y#]���� ݁z�7��u�8:E���@��c7 �i�wW����qe��|Ѓ<#!ݶ�i�Li9�'/"��C��,`jj���x=g��4C$���-�b��'F�4�K����ȳ����pr鰹�O��9 ��#�7������v�R8��6j��|�,σ�1��9M��Y:�}��6�ټ�oY�4!����|[��wOp��1��M<zX�p��	�w���kO}u�_��N��;?*C�p��͙�ۺS9�HC������c�L�Q#�� -�QO_�hnu�1�_��W�9dO��On���Xx8��rP�
���"�č�蕓WTr<C��>�1Y�#�_��1b;\!��p��EC��(���uy��غ@���=���_҉ݦ/\%�gz��X�
ٌ`7^� ?��B|�U�z�$����������bB)Q~��EY�^�;a��4�~�nm�ɺw��<Z��=NX�Ƞ3�H����B��[�H�;)u���l�\���!ɑ_�
��%��Ɓ"���$6�Ҹ�b�Z6�r�*�5��UQY����6��aL��+��v��<Ak܏�8�GK��m8*��a�HD��{��f�
݊^s"7�����r���oV	�q�!k��'x�9��h:<�e�*ft��U�n)� [�*3��Oύa���]k.b���+�}8�  s[GB�R����|W����k�M/����K:�i���{�fO׾�ıo5Ǉ Cf�[mU^o��6�e�;�>B�L��oԎ{�J��i�A�t��ͦ$MM�2���O[(z�w�W#V��X�Ѩ	���3��`�g��e@��ͷ)�h�+�1?�_t)큨�sƜ\��5Ͳ�v"ǐ���aU}{��t���z� Jo�E	(5�fI��W��b�zV ٸh�%�o����?��bG��W3��/[�v��2L��V��B\I+g�m����){2Ew���w���G|�$��T0M�e����B��IwL�_N�ta�Ç�|{
�a�q*1]Bqv�,M�x�"R�>Eo���Y��>�!��LZ����u9!|����܏*~̾��l}Z*�����o]>�6Qqko������A����r����5esp��P�A%������y>�fIu�f��N	�ӥij�*�W}�G=��PD�zR�q}wM�ʢ���V?@��g�\�Hx���^�ʦl�m��q5.ʪ:2�$4�%�Ub�7�0��|"��D�FSD��dq6)�ڒ9��PlsțE����� n�$]c{먢Ka�Feb��M�-�����T�{������dn7��m3o�8dsЙ����x���f��n{~8���c�W��Xv��)����k�x��^�&���W�R� Wھ��G%�E ��֋j�,����!P�<��D�M�B$Ӎ�ܫ�oOY�%������9m�'Z��׍����C�����.�uCJ�,�Jt�\QDgM�dw������3򭴹^�_��q*"ym A�im)ݲM˵s'����*D�x,5E_���L�.Fv�4/��>�D#=��H��Fߔz�ߓ��_BG�&��xƕh4�v�|��dD� D	�>D=�)�}�h�P���Ņ%��� �\������5!jW����9&Q�yw&��F:�t�z�5�T���"�~��rr������ޱ�О��!��E����k�/iżC{��K��*go׫#����-ϖ&_E%J�/���-'z��p���C$m$��x;�1P@f��>7ĸ3�o%
��ð����A6�%᷼�]���S��߇&X�T"��)��ۯ[�'jB�0�z(.���t)�iqz,�B�ŔeT"{"�^�?�&|-�+�Ka� b�	"zhdWōн��L���t����t볡- (�Y�-t�!{���	�s����G��]F27z����y�� 9�	OD`5ʦ&h�!���d�X�!�VPuh�~uď�c�(�|��:���8?[�~9�JZ�k�kW�Y�,��Wq��w�Z�
伊�By��6l���Hz�����*��*w���(J�YB�.,X�n*=42����z�1�ω�;ܤ6	�uA�ᭃ���8G�<
����@�K����om����8(�P�d�%���~�@]�Ds��h4Ƭ�������fא��.�
��*�uN�U��{^��	*�.�K�|wrD*O0:��I����"Y����C""%�!Ԋ��yB�w��xY���4<��r�E�b7������3�<�_��g"���'�i�ɏ�&B�"��P,Í�(6�ΌA})9�����ֺ֘�՜��t 

���x-ױ��B4��/�jUOD$��XD��Id&9�������e:ԫR2ӟ�ZZ����p/7E��`�05��ڠt�oW��8�{�
��g�[����	�Gn��3�)�?z��?��T��0g"�_E:R�ؽ���FD���*��1�?��t)M�|�T�BM]0k��*����D$`;,�c��NB�X#����m��rщ�e�aZ�u�3W�-��$��ƭ{�`��
JБ%Q6���$Bu�W�\��E(�2��C��MJ���X; ;���D3GOR���X�����2�S �[=��8�*��x���'b^�T�鋠�}�ʀ����m�Q�2%��9ZWt��U��;��N��l�2�*�-J~(������t���.J]`���= N���'�I��Xf��9Nr���=N�n � � �e(.y4��k�E۳�W���"�[�߁��GH��Bw�\�X���b�o��w�r;�Mi+O��x�<�"����c�J��gc$��J�5�حW}_X4�!��.yDC�|���x��&4VtB�R6z�k����AՔR��<j��Kj�	��S/P�����"'�pV������S��Q1JTB�e���L��I�{������[Ӗ߅��'s{t
jV�8꥙Yaxp�9���R9��[�Jϋ,y,з`oY�PJ���0[�W.hc�����Lc>9���M.J`����L|&��u��u><�JJ�����P�^���hN�^���f-�w���Ur0]3�t0��������𧇛aa[�`m�f���	���:h�y�e�Rq�)t��חB��u.?.C�I%��Gu��uk�� �|��:�4�\���4Qs:�!��n����^�w��D��=}y�So~c3�*� ���ԕ�U���4�c�R�}�A��`X��r�,C��c`Ј��㠁��(��]�g��3����3���)�L/�����I%D%��O�Q�J���Pc´�,_�fFZs�3����'L�"9���O%v}p$~[��0�����O2������v�;�����7"ìMǨz�����e�,t������-�F4����T%X�ͧ�:��I�P?�H�O	��*���Q?�%V�O��3�P��h�`p�9�
L��4U��,�2m=��M�o�·�E�c>�ɒ�dz
�E�>M����S�NP�s�pXM��Lj�^�Ƿ�MC
�7W{ܸԕ^��������WI���lZ�����|�8�f�5pCA����a�_�������ԝR����}P��GP��D�t�s�v���Mo�9Ti�A��޼A@�\rؘ���G���l^�)����"B��{M���~\���R�-Q���|��%Z����Cܨ�r_Z������,�P=��������i�N@�J�=��n@ 79�� ���s��^!]9X<'x򓏄&a����&�n��j�ז������#=�_��<���|�_^�r�Hb{m�3WI�G�v�[a��EO.U?d�S^p�&�
hQ�|5�q�]<����YƊ�1��֖��664����,������J�&]e(�=�Ft�\'Ⱥ_x��ɧ���bME�g|��0��t����
�x��V�J����ԷpΒN�Th��)W/������S��p��U�BL��^�U}�NFr��dFId}K7��F6��nGG�Ϳr+�}�\�T�7k��Um1�k!ٯh��˯�֦a�P��:�������L
nk���pٯ�	�E+���?k��ҭ�k8\j�25N�e���(�n�E�w�{]���3Xꇎ�6�k����Ne����m�4+&��|j]�n0VT��9mТ}РmNB9���i���u�du"Tn�>�
6�)�8d��B��0�Z�X���8�ܱ鼭�0XS��w��)f~����Y/���.,�?�*7�c��VS;��Y]5B�'��M�J��N�2B��/���_5�;Rhgז7mf�HP5ܐ�"���%5>�y��`<$O9	�`�(B�+�T�:xt���8�����_p۠��%�}$�\=��ʐ�:k�	��|E�=�(�I�d��ĥH���N����?�)�v����7�����ۦ�0�D�@8��Vd����	�'/Z�e���$�ef&B<��{��k`�Yaw���a�$t�c�hs+UR.�Hmm����R!��Y(L�X!��/,h��Ǘ���̓u�k"��U��[epә�Re�(��PN�B�b���T�_"����T�DA�Y�y������F`z���B�)	^���ݗU"��d�Y難B��J��&��	+����s�:HC�V ��;����D5�&���Wp$� :Z'nl��7�:rl4�-Y��ш и��<��%1)o��"m\Wo�OJ{�Wt��]8�Cv���XP��m��m��8�E�:��lr|��7k��gc�rfe�{�M���B\�$�~��eϯ8�Ր�M�	@�	ʏ�=;��\	�I�M'yaR��3�
���k	��^e��f��h����Β<P���?����FĂ�a�L�z�K���7+2ן�Tk=-��+�ޥ"�@�ِ#%쐳2��n #���
��
a��y��"N{�sS�YMu�ڢKl7��f��D��;�ǃ��zi�~��3Ҝ0�\�H��ZU|on�s�;K�z�$��]�q�����T�U��a�!�<��aS.Pj�����L㉴U�� ���	Ɏ+L��P�����{�c��z��~P;���j@sWm|�������$��ZȢcC�4�/*[�-��o*�0�w`��Hb��f����5ѐ��\�Q�Qp��򋨵2�yņ�	Qu�c#~ﵭ>���vJ�>l��4��� �R*Fr"S%��ԈZ��GEJđK5���1��l���n#N����\
Q*b�0�֛֋�S8�=�F��c��g��7���CV�|����<�B���XeXr4�,d���7�g�q����J,wB�G�[;�61�J7�����:�@/����p�8,Kp�y]2�x�,�]�������|E}Lw��s��S���4.����$kU�d�P���2ǣG�^��;HV/-�7��8V�s�[~��L�`�3V�!��P'�r.�D�i����%~k-#�������_�@$cC�9�~��Q�rO۴Tx�3i�|
B��xY�ۖ�'5�m;0ӈ_*W�.��<D;jE���ۑ�Q
���P��YP�B3���]�WadD��UO�� ��2')��'��bSr�v�c�!�+�
^��e�\[�w���5�W<������^���C�-���[�5U���專W�^h�&T

b���[~\x�-��<�3$��N��R�E�f�M3�h؆��J�`mi�Ϥ�w3ү_|��iˢ���l�閥ɠb��[(��v� ��v@�1&���g7c¸�<^�x肐�
\���C�oc� I��~8��y�c,��'c��|_���-1���	�gGI�Fy���R��w_t�R����9���Nfz)ܝ��$c�Z�I�&q�]�j�!K�E���;�5��	-�����[ɲ�%w�x}W��눡 /(�?�m�,F?Yr���	����W?ۭ�SHͦ���3:A!O��7�}QN�8�N�#U?])��.��>(���K��[�����:�'�OD�6�n��� /:�@���k�@b���Y}�3�G�n�/�q���&G�枉D�?��E��}�y"$�x�n��*I�pz�, �:>�Nv�TS�+Z�δe�]\��_����7Z���&>���F��p-��b��T�8�t�}�w�����R�q���Kȋ�G�P�,g�k7ԝ�V� 0~o���[e��c����	���@��6%�Q�@;�郮����D�\i1D��YL�=�/G��)%�����Pg�W�O�>->T"l�QXO"^[NM/R���AL�B��a�E�]�a��
����z�	���[�����:*_t�_b��ܒ�x�D�Z�zb/Sk��: KA#� ˅-N�x�����������m��#暠K�8$R���f}0�Z��j%&��԰�
1�����G��2B��R���]�@�?%g�u)�/��;��PQ�xM���[@}>�x���������K��#��,� H���#L[���� �S-u��9����M7NhCnYpc~`g2y@�eGs3�I6���̠ u��u�$�\�;�9��e��`����,!6��ˑQ}:�lL�o�\T���� "���o�Wc�>�d\\A��Q���\��� :h�ga�90U��'x�9�`��vJS�i��$��W �R�����>�OW0���Lc9m�����xt�X����&-��\3Zα���p�6G@$���R��+A���{f�<Ӯ��:�*���ƖPU�`씘�&!���bp�(��+�ɸ&\G���Ia��>V�O�����W��u�_�����'C�He0���?y�W�/�5�R7�9��.��)�j`���E���,�#�n����yv`N�� �=i(�X��#e�\�q��P�۱�ғ�^�w��.i� ��-Fo^��R�\}}5��&8����;�k&wuPA�ViK��[z:E h�Om��5��1#��;,�3U�����4SMADH/ ���id�|ZX��>ta�x�[��?(�$��;fD��K.�=ka� B�ɘ
��`��Em*��x�Юf}�2s��>���V̓��Y��!�yǸ�ʍ�"z������ID��ģ��aa[�8C�'�x�Z�����y��T�]� �aB�|���A���V���PP��x|�3=��:'�8�<�\)�~��z̙qf�`�M�� ��6��E,���6���-��|)]tض��]ӀJ�L�߫�hR�Y�D���S�fʷ,V� iI��z��Q|6;z��vY%(Kp����&��L�#`����߲ؽ��{4D�ecM[��\3���?�&�2.3LO�@��upgci���m��*=��%�/n7�!ϯ����9�����;Ԑ��L-2�z��ٿ@6�]�����+?�{�"����r��1]=LH'mp,(6�qs����͋�(7~5_���=+�0��Ҩ'�H�s���m���6��QO�&rV{4��V�Nt�i��;S@������lz˪ナX�A`��T�V}V��q*GѮ��d�\꜅����zv�N���e�	��Τ�[��X4�(rt˝�G�0Շ��v�n������R9�B�NN�몎����E��K���Ђz�H�FN
�����ZSM<jb�}��k���_��ݑM劌c���Xݟe��?�^�)¾ow5c�c��d� q0n�?.>��W�+:�{%}�r�$�L~U��f⌰N���hmJ}|`Ln�*K\�Ή��V%��BVUH�ua??���lZ��&�
�/W�&\A�����,�6jI(&&�!ГE��.�J�!��v�ഹ �N��\�0�k�X���Wǜ��d���H3��\�$\[)��:��k��_������0|{c�}�r��Ar,B�C�q�z
dp[
�Ɉ������;������c����>�-�ok[?6x��7P<(��)ǰ��O��t�N�`b�#���z��V�8T��1j������i�w?s)�	�%��A;C�1Hφ�сii��?c&��esT�a�$���`B��ٮy{��?�H��'!���)��,��l�>��Υx`���������Qҿ~��a�
����K�ZM�%t�*|���5%[��%�䲚�ꆺ�z�'�c���_ʒ�i���^��<�'.�����:l4e�,`��7�ZwS.*���if��T�����O8�"8cZ�{$�}P����r~V�Uh�l��k�DEp@�Xzø�h=�>���F4���䑂��Z�2�dM��~�M��:�D��ƨ����33�s��L<�y\������Ui?����>(Л�2��Ԭ
01RdeY#��&�DA������o/�3�?	���/���#~M�Q����a�Н¬+SP����6l�	����J4�k~��.�۱m��@�fq/g��E�����2�9��L�o��_/�'��c6;lMvT�w��5��$q� Y
3�e���� (�Fۄ=��i+o�;j�ɾ�>77��G��}�S�QE*�Rc+x�*��&D~n��� ��:l�!�����"�ʹ�	����F�M���8n�^tt��r��^gQ�	�4h� �ٔ�ܰ��\#Q�9�����@zA��ћ�����+Q,n%G�[��`����zjf3^�J��^˜V>~�;��O׆��!Ԩ�� y��E�
�/|.|�-�"��n��%�/�*5wg�47���u{��L��]����DA��/��H��o���܍g7j,%�}.x�N�0Y�ZBb�c17'�6�/��f�~(�w�s�_݀0���mmXS��̶}M�[�@��~h����Zz���}c�m��x�����:e	�����k�pi0#�b��[��u�����m�;H&���*�(R�c�z��X����ʐ�ئ�bl�k��ɧ~cdiX�
�V�0�Bb�;��PRi���Q/�L��}7ߐ�'.���C�z#w>T+x�K1y�"�y��G$h=�>P���r��L�`$��0��p�x�4hQ&7n$	�uPŐz*�߲��Jلjs��f4��~ۓ����\�
t�/�Tt��؈�>��܏�uV��M��d��H�'�"&9實K�ʰ����n��b=ط`~���c�A	)r��� �PO�ʔetUq�F�.�j"�J*�ىꦧ>yf��C�w�M@�y:�������I�wOh[rا0ir6�J���8�<�+�?BWq�ш����Ơ���E+HD����QS)3qf�*������7�[1^��I$��/��|}��:����l��@ir%Y�(����s�[�R%�[��u�
qe�r�xD+��`ģ8�}S�̸َ�ۇ�Ȧ�C�5�dO���h�u��W�9�Ml�[�g�ղ��KFl��r>�.`x�&���іXm���%<�e �(u����^�B�>��H���ȯC�ɖ�.����A.ۥ��U�V��~eY����wE)�J�7���A1�Q�.��#��ʭ"Ev_1�Y(���,	Ŗ�.�	�<A�[�ٳ��hCn�V�b׵�(AQч֣��?|W���ƕM�L'Q���y>L?`�"���������6��Aېt�=~�p�xg4�5�=�+P�ɸS�j�zuD���//��dv;��D)�IX���ۯC��H�x!j)މ͗���N��|Vb�g�%-�8���$B�S'�)�a����Ӆi4�3�Eߋ�煾��r�F����cj��ȉ�.���NH�Cp쫳<�[>�#���m����;-&/�)-�pä|_}R8�r�C��u���k�����f,���i�y#����Bk����]ܗ������$�G��)d��dT��Lt���@��+����3�ʒ�#S̣��KX�A*�&��u�ۅ#�ZN�\D�>9�jB1���Yv�le�������l��V�M<BBj+^p#�V&d�ɞX�n͠��O��a}�%�i��W\Yva�q��~���J�]����Em B���/g�+��q�f�<p�K�QD"�>"��>�c`�bLl��W5�,rV��[]��2�t_�3W�̏�-��;�6{�B*_���n<Ðȟy���|�����ً�d1]��x�]h���`��]��޵��gh�WR!'�H�:0��o��i"a�*�>P�8�#�� ��A��K��
�E�թW^���SSip
��w��{���t���>�e��:7aw�Jp2h|�U�>J[��-�(�a�%�0?�K�|C甘KI\:.��M�U��ɪ���;�&����������}�b�>��1~brN6��釢m#B�h���y�x���7t��f���|���,�CBᚅ5 �P�3�]����@�@iH�-�K�y -�S'�2��F?t������1�S�L��� ����a��Qԛ����9�d�̕Ś�$�4��ܵĪ^�P��=�pzl-�]�'{!��2����S�@�S�A�W�\/�b��q���*�&�^c�/q�Y^��%Vp�&�2.�3���~�F]���fT�!;cP#�t�Vi��w!�+w����SS�@���a]J�Ձ*|��U�F����ά��'-ͨ�6��d^/���6��h�ԭuxTX\&7]x��k��~6v�w��pF��m�9ܲ����%���<Tf��\;IG<�>��]Uǻ�V�S�u6VS�D�$_��t�����!�y�u�ޑP��ct�:v2*�5 �~��i�g4ꩁ����L;��$��ɵ�N5ޖ�#���s[���Q� �.��.f�0$x"�����*Vg��B�s���b$}�3$oi����4q�ۚ�V fr�~ �9x-L�Hs� �4�љ�����<��r��",H�9K j�Y�h�G��.�.�噲i���b̵�A�h)lO��R�O�BRzyrR���L���*�����?���N����?B�����Ye���I6��3�d(�|X�9+H������1q�|i�x�]������Z/)�\��(�\L��sR���]�9e�M<��������΅�l���^�o=^�"ag�\L U�v�?h����NjL��W���>��?�uE�V=9l����ǈWR���;)�b)g���,���B��t&�QG/����9	�i�����hA�	9���2-�����b��>�Ï����R�M�W�Ʃ��:�����4e�(��X�e"R|w��C���]�QU���:'�r�Z��QVq.�C;jןP��]���>5������g1���%��+ܝ�r�ЯX�>�T�9��f���G0�J:�o������-]��^�p��,��:�H�����F��Ku1��AyHn�v+\݅�L�ZwD]���n�=?xLpU0��T��hZ%q�]�5�͘=��l��l�y����l '�б�5��yغn�B�?�A�Llx�"Պ��,��)��5)�U91&T"9ɵ<P���/ T�%E&5�#��-��/��;�-�o���S����u&�Yo�骄�5�:|5�\�Td��bL�y=���^��{Xu�����B�޷��������2�w�B�}��
�0�M���(C鱣�ؾ��8�f���l{L��W�M)3ѩ�P�a������l��̈́�=�5�����#�ZgR��Sr��&3�O��*���#�K�G=�O��y �+ge�դ&8E*��8���O�M����������rxp�B�B����_�w8H.Y�eM.0=��P^�=��{h3N���V�2J_!^_?�j�eUi
kS��i�^�ftjA	+	FC+W�Q|C`�0&�Q3Kݥ����Fw�������Q5�{َ�h,�w��Z#�[A�sݞ!�T$IO5��)�K�
:�#�?���laeZ��8�Z!�1�o�������f���[���VQ{p�*ꁧ����YɵCS�V���[�����K{P4�����]z�L-����g�[��Ա?� ��ջ�+M__��8>ȼҢ�w��v;n�/�S�{�� ��y�o��1QKs~��Z��;ǯ��D.Ĳ��v-�
t�(d�O�l>�'+f��ΐ�~�%B�zI�1�xo�p��#�sZ�"��g;������K�yo�M�i��?���&@�P:�˽2�O�a�خ'֑�kÀ�}������Z�dQ��cE�]"�ԥLf5)I��sMx�TB�4h$�,��f�����t��3o���Fy��]�C��'_ �}-H�r����uؙ`�#U�ڍS%�1j_�y5�2����*p�iҭ�����r]Q�4�x({�)z���0�G#��-�X*��x'�2w`��?���G����{�=d�7/Q��;�v[��Pk�е	�o�)$cz�($_�"�T6=ѽ��a�A���$ऀ�-)���@�|Um�t^>$�uwy���ч4��9q��͌m�ߙq4	����í��q�(�	1�m|�Y�k|ݸ�L�"�<�h�|�	��]��M�s,��Ҝo=ɡ��H��H5(!:���1tk?�6��c��N?�9�5����uk�r���`��i	M�lk� ��X��y�,4� 1���*��F�3f�K��F(Y�
�5qV7-��v� ���b���{!�g��,�ݰ�ʌ�~��gw�\z�g�`xFk���_�>�_����Vv5?I�����s/�����xdtpP^ףּ�Ӷ��ld>�:Lᚾ�	L0C�� �'�V@5���WAꤷ�y���U�a��� �J}���IN3J�\����J�,C�ᘑ[ٴ�H#ѫo��̍�	���!�L�7 ,/csYL$ ^AusW��[%�Va�GHB,�aq�8�a<nc�e��,��<x�i��oU��H��O_�/1��$��ހ�A:S����ٞ} �#ջ0���"��wB��*���dnվ�lg�.{�>��2ѭpC�	z�ꃊ�����n����w�
6s��#��ʄ����]v���U�@�yg��P�k�]٬�o�2�G�q,:�%מkV�tyJ��e�Ly٩t���X:�����g�*���Z����j�J��r�=��[[�YI�A&�~�a�D��AF�m�N��o �M�Ug�׀;����/=�ps��D3�]�j���Be�!�/��)�K~�V<.wc`�ՀFC��X�FF�>�c62r`8/�I���O9�7��~q����S\{���p�S���Q��9��R���oŴ���UB�ƅ��ђG4T0��M ����a�N�9�k����T��,o��D�j�@�X�����K��o.�n��]u�T�Y'�iQ�-n�&����$����(m���IG�H[�10�.����l�p��xz��5���z�TL��1���?^��8��+u� Ob	=�MdM{���4�O�*������о
�S��3!6ޔ���u����[�&��T ��>�n�B��Rϼő��[@�䘔2XB��~4���1���\�! 8�"gc���{�޺��n�'��DԮ���U偟�?��:z���?{'�^C�Y��T%�̭��%Kp��h=�(B1�M7�#;$��QZ����Q�l��g2�=<���'Et¢eZR�j@v���Y¹r2�B1A��@��n��[��)6�����X�=���LbG>��1?���}:c��l��8
ы�N���%q�.���nÆ�'�>�4鍄i�$o�Y�ֈo����,���&�Rb�D��׸�b�N�5�i��ᨓ��,���J��_*��ud}1��_N��1�!�AЄ��i����\�Z��L+)�������L���JUb
���8o�)�a�s!u*{F�̯�4�#^�(�{.�EGj%D�&]69La�̅��-{��m!Iޭ�!
8T��r��8ȶ�i�芬��-	�|C���+ԃ��z�w"Iޞ5䉲�m�Z�l�G����5���GM��XNv�Z~��Lų�g�`�h��J�;�C�@*�� ���=$�X���^�X��rA�������� �����5sb���`2ͫg2���_�~vHfh0[���k�G$�D�:7�jP?��n=|�Ko3�~�]��]8#����J$�$�M�S<S�؆9�#F�'���Q1B�u<���h��Q� �6�`��9������yB��[V	��)�4z��%O�7����� �x- Q��y���T��Z�݌���0�5Gxc�Z@�]�$�2��PQ�>��{2xR����٦w2P,o5��H��0�r;-�9*����=W-�hz�==�Q�i �QmD�	,H���ʥ����b ݭ������.�A��U����)�&Gx#=��/��Ě�yf��h�Pv�d^��D1��XZ�N��c/m�,H�	�yd�,��^�������x�(f3F�J�Y�Rj����k/a��t8�VZh����fk+2�j��w
�r�e��Vspޣ��QFW\�݀��sPSyT6 �<"TP��y���ee ǿ�>C����U����))��3��`�`<��$�Uǰ��_X����Q���5bt�7�Az��:'�T��^6 c����x:|]��s�H�����:�<,i�X�Z��v�K�d���l��|yB���$`�~uB&]�T�s�O&�fE����C1�̜���>�Z�ju�%r�W'��sȝW=0V�[-���eb��
 ����,O��$TCMz��Q%���V���Ϥ����\��PjM��CH������*�!��a�9Aw̩���t&G!]��>"�pl��K8b�HY�'��@�U�Z�_�`H�|�f�L�@���l9|��Qsd�|4VjY���s����I��%�7���O������U�� ��dSvFԅ8a&��0�3L����T�eG&t{�2Q��`���'�sLLf�<Uz�
�C��/�F���ĝ�r�ꏹu�V��l��N����M�0�{��=pTr�����,�ÍPxg���P�2��(��k�g<K[Z3�����s�w��W�;nR�{Э������K�e�B� �,/���g�ʂ�oø����IG����{ǥ�N穻��F���|��0?�i�˛��-֙́�qT)ծ�}{~%�@B�X�8�nj�*u�<]�\��F�ݰӥ}�OmwD&�>Zԯ�/83z���<h��=���e�k��	qо'"���ė�����
�9aGgB�����h�o����R���Rt�̥�b`7�<V]	����o�Ma��tݠ����G����h�4�r����Ȏ��/%�p�+#j���O����\Hb��j
���u��)��i�
�Gj��e�F�$Do���O:`��w�Y������u�#�aM��jY���Y����<*K�%��\vޢ6�;7?�Af�Ć��r�o��Nf͑SX ��{�ԕ|t��%�̙��m2�Y�_��M_
�+s�yH�s`�S0�	&�Oe-[Z}$�x/�x��\$����6v���p�Z�w3U�l�!v"�I��2˵SYuߎ,�>��?��&T�jq�����b��7ϓ�#ˀ!�5��k?��s+H^�9D��]����bWPU�8����)��C׎��D�1��)�:���ى�8�'ɏ�a�o���h�e�0E�;7!��z�sWv��-���9=��hїV�T���5��X#h���/�7��_Ak	�`��T4�4����!��nm_v_2źt�i{���DZ�X�Fhgdiߡ�!���v����Iy���������Q��8�d|��ׇ�zM��\�J���Yp��(ɁaG�1ͱ>U�
+��	A�@���ޢS�V��K瓁؎|����Ay*��w{�j��fr�2ְ2��ݝſKw����U�}y,�ȕ.�*"��"���if����Y�$`��5�����1�FfCD9�2~����m�X��������|�#:�IEi��0��|
��L[~i�=`/���n.+GH}]'��g+�b^"�:�w��Z�Ay���.P&�Ӌ�
O�.�����l6���S�&��=�xy�ph$0�$�O0�W��:4oU0��JP��'p�24���t�7���?��P�.+'5H����9����z7dw��y�;aaע�¦������0��Ps;x]����a�+���-m>�ZP�����4�E���-\0��֘��}��L���4���
nu1�yͤ9��u�()LXm�Ẁ����r$G{�7�ۈp��Y`���m�j(ڄ�����o0�
5W]ם!�7�뛿^ߝ���_�a b�}.���n?��Hu].��΢5��-d7�c.c���z/F^�ϐ)�Bv�	�zj䷕ik��a�qWtb�Q� .9KkE����n�%���=��y�����D�T�%�w�5��w
d嘽C����&2����*�.);t���sH��j����¶����ny#B����:?ԃ��P�Q�TG<�KfkB��&�haP,	����ݜ)�4�a�"8A��Ԗ�w� �,�QR`�0��� K�	(v{���\���)�[������v�8dX�(�C���/����Qbe��#Wg�K9M�����E@�@JK���Oڮs^��v(����p'��n�x�:�kER/��0��{n8CU�I�)�)a>�KNϳ�������Y��*A3���Y�k(K;��ZJnI,y�g�#QF�L����B�kQ`�l_��6ܨ>8��[�$ȂOr�[����Ozx-�?�K7��)4�{RBYy�%g�}�M�n�J}X� �-iĘ^L歵��e�`�t�)z�rQǹat�g���m�}mTM�T��{V���h(�=����rY?yc]��r�g,.��W�\=��)	�*�&���zaq����}�g��AS�cv$�P����j�߽�mGޕ�̬���M�i/Tx��Q֮�q׍�����g/��>��4GZ��AC��eM�X�������VC���~@����$��f	�4rK���2�Z��-#���j;��a�!/�! �SM�c���Qm��E�&�]�҆�=��YR�A}ֻm|��,vQGOZ{E�	"H�B,n���[)c�<����@��G�jy�f��jH4.�ѪRS�MG��h��^��n�1sv4Y�v�UC0�͏K��M1�kc���_�����Q� !
4�&��٭P��{��^B���a1��0��0�vy�r�ׂ���Ɂ��Ū-����k��>��4����]=�)�b�|+��F+�d�ɋBG�9�t+�(?2W�@��7Q
���0��q�B��q��Ϡ���TK��GIѭ&���	�Y���wvB�"،1��ֽ�SfET1�w鎮y�(U�eXiW?��C�v��[2�I2a�&��$;��m��f��n�r�K>Q
F��CH֕� P��K���Y$e].NE-����΀��`TL�|a����Sz�����9���xë+���p��jq����Hq��M4��[����{6�5�ܠl%����^9�b}�<H��V� ��أa�4��������'.�%���j�[.�Ȋ!��)�+��J�^R�Tl�r/e��7)`�h*��Ϡ��GDB�d�D�bԫF�0^�b��󵛒�}�Yn����U���B����%����bx��;�l�b�e=Ź�S�Yc<3[�A\�Rݻ~��1���8�Ā8Ձ+d����_AWN�U� �	:YǣM}p��@�^3�*�@��P޴�q���*W^��2��l�~]�x���#ޯ`U�V�k���䒏c&���l�GigbӎX�;��3W��sCc����B{/���x�l�����h�j�t��W������>r � �'WY"��Wj<Q����@���U���1��h<�q��/f���g�y#���VQ���7����l�=���X��1.�\OXp$����  �~5�b"(�'С��$:�X��1���o�-5YN��ô��Z��#���7551��qs(� �̃i�omѬCl� b|>���ȚJ��d_޽Z��^B��r'sڍ�����a_FO�.��i�ܺ�V�|�������ѡ��SI���
�|M>�b��Hxe�6���}���z�|8��s�������SV�%��:"���C�В��	��8���y��en��Ex@@O�B��z��
�I�%�LV�pDA>�>��3�3U0���M�؉�NlMޣ!��ҋ䙄J�B�R�@�n-}��Z��"f��:ck��S�"U9ʓ�J�Ʒ�*�[���8��̈́H>X�k��!�",]l,q�6��7z�R��J�) �S�إɾ����7y���6������i�Y�B���x�&���r��G"K~n׉��X��Y)y:(��-/�˝�@hQ��Ճ*��-({��b���C�����`}Ì|Qb��c�-�����#�m"��u�#l�Ve��u"fl]7��ʎ�]s�%�M۬h3x���P/w����-8UM��?�To$ZrsQH��C<��!���q'�_��y�}Љ\F0�)

��ְ̀�1j��[�\p}%ϟ$T�+͠���[��q!�h���x"�����r��7��AE���' �ڃ�a��Qo�����'�c���F��;�س�L�R(O��A�ck�B����3�5��y�a�j�R<}�1�y����s-M�����NBK�I�ZV;=�~WO���K�-*e��2/��f����s��q!���nrsOCX6�L�� ���*z6��1��`I�G)GI����5�a{Y�=�E���`�����YV��J�T��^R�(�;>��;�9uV��.v.*k/�r��8�w�/%⏜�V&���"���U�������ȗG�V!]ޣ��5ô>R;��A�����e 8]����g݅NTӵ�^Q���~G���@�k���<3�d�=�{U����Q�/##�VRpD{A�%��
�;<���g�.�Bc� �k�(`ш ���*,"T倈狊Lr*Ć�U:�Z �,�e>����P���tqNF��Gog�aKgOgH3C ���x�Aq�$�X��5�/�<����j瑪� =����g�2^5H	�{?.��^�ۺ��RK:��8�jzM���n��� S -܇R0�xҢg�C�R��!o��­�����x�֡��s�x�Jɉx�Ko��1���*��G�]��h}�V-T�����$r���@�V(�	9����@�,1E���������Y�v��+7Ӟ������F��ne�鳿I.b(N!�s����+����ݔ����JV2�Ʋo��<��0�U��1���`��=+B5sC��Ig��� ��@/�D"DjP���#$�����'��p%��\�_w��8R8�1~�JC�=�_��~� �Ё ��k�T^�	�^��ƚ��A]iXK��ٷ���9���n4��<4@U��n��!_��*�
&E�Ȗϒ	����uy�id[j��  a�8�^�}�U4�P�N!�ip .�u����m�$�����Z�S��,"*��8[���Η���1a�ghJ'x,G0����eM���ytRa&^W��y�[(�{�Y�s��5��(���*���.���qV�}��8��
�p���Kڕ�B�z��]��jb�L�e��D�̰\���o�N�`��=r�>��(dE���HM��^����y`���r�ޭ���~��=��ل������+��V(�b�qyb^����(-Qʤ�T.P(Q^ދ�#�O�;�p�֍CC�G�(F��7���1���~����!����U*P��<����wi��Y�hb�3��wL(`�T(ڞx�tE�d��{��m����0��+Tm�6:�ݕ��������^J�ɉo�^1}1��:퉱� w�^�Ȥ�R#z$`%���/���ؠ�����ru�q�t`@���kC��B�op��`|ܜ������u`[-�d(�p��b����u��Zzg4oͤ��DT�@M�9�)"SBK;��s�h�O�@��]�JLȫ
kau������������Cg�Sod�r��ⲑ�+XNјF���X�;�]w�	��p�TG���P0Ew~��<�}ƏȈ^���8Wz	��'u�5�ܮp�x�� vL=F�3r��{~�>�d��o�P�m��+�:�ح��v�Nŋ���"���׌���0�Pnu�k��� >����� r:u��oN%$ɬ�<�[@�o�X��Z܄	�'����n��(k�hwT�O�E|d{�H�؇�<��C��WB��o�͋+�����ϰ�^�J䰦�0;a��Դ?pk���w�h=��;w'm��;<4w`��We����R_�1,@�3f�@���@Iv�)��i��P�[a�'L$|�A_<���'�bU�w�B<����P�ÞD��@� *F��{�4�j�s �GD"�d͛,�8cv��8W9��:�'*
Y]Z�1�G�}��Sy̸��q����/
eC������p�4����d��`���<4�?���,,OC��)7Vǋ��u�؈LŎ�P�0�� �ކ���w^��lHR�'�D=��������Ы�=MP�� �'-��9e�e{�����4���Gm�yqB%mn���x1Я4j�^�Ćk��q�$^��@s������1V������Sƅ�c8J8���@�0����A�q�1�	�FC/_S�j��C�������Wu�~ܷJڻ�p!n�|�}� -4u�8D�	�:��8�#��R���{��,��]	�W���5[L�����7�2�"K����P)��fi��߹����&��V�M v�\
e�TM|&�ɸq���!��&�f���߾�4�����C2�"�4(Ċ'Ue[�y�icwK�t.G�ay/�I���Sc_B6ULq�ZI��QTy�T?���� 1k�; 2'&�� �Ӟ��������}���}󺈞wc<zK�!��Z�Jfd��#Hp��"xa�3��,�Fzߕ=�����
y����}b�kq���8�Y���f���ǆ �]�vE��%%Qʡu�v�U����N
�b���N��u�j�$ٙ�������$T_JX�\�z8O�Piªd�Q0�m���Ⱦ�[/|�4W�a�'�����n���WǊ�t`� �h��"��NmQ�#ˑ.��
S��{`Hp��R&�מN ��GR��I�4��a����(w\ĳ�v���c&����:�orۯ",���,hrQ_�1�wrG�a�7%�YFMZ(&����}a]�W������d�S�=)�.+�ONx� �HF�Qr���*j�����@�(���EV�i��t4�����r4%n�Tc:㔎Tՙj���_8��rJtcXǅ�8�C?��&��1_-2��P*"�9<�I)c/0]ܠ���Y�Tm�;�ߦL���Z��7�o���6�������N�ӱvn��n�TV ��6J*Un�~�٧}\Ո�V�v��㿖Ţ�ѷV�Jt��y�@����|/��Ѷ3������9��E4Q�vէ̌&�����M�jP���J�`�&"����*՚�����~>g�H�P'��X��/�L��H�'n�5hrj�B�U7��}������d���V�J���2��f�	e;�nH�*Ǖx��O$��ݔ�?&K'|��S�XR��*d2O�$ԯaIj̻����=A؊�uJ�ť�֌�)��	r�Z{0��j^7��e���3:�2��0��2��èL��]ֶ�+��F�������W���i_c`�,|�JI�T����v�Y��"�J��]r;�t/�=%@��.��S�Mt�<�a�}R��7���X`��B4������_�n�K+�ˤ@1 ��a��˩3'{�C9vW���;R�o?H�K�s���j����t>�|��Ua�z_�W�Ѳ:�C��$���e!;kv4����.�����dxa����;�nAs�P�����F?����?�m��oj�����Ἕ��T����f㴐(1��������G_�(O��nz�1�~���#�%/�{I��5t�r��bp�M��C*\�6�@ĕ	�/6tcA���7܆���p3����Z�#>%��C��(t��d�2��9�A�A�Ԍ)ڇx�(���9�����$┛�Me�s�D�r�[������%{F�fۇ�z�޵5�$��i���RR�f��T����Զ^�|�H�a���{zr{��Y��^�I� $��婧B����w�4�n�����d_4��r!�F�,x��͔�N�a,����a�!���f�
�����q�EIp�dn�Z�6�ZN{�S-���h���҇я|IW�u���{a9�gg��M����a�M�f�̏ ���_�v�s�%u[[���ϻ3���L����.��a�(�p�m�\���V�:��,�r�)��4����^�Fve\7'�9�	}��Ҭ���ף��U�,)4.�3}B���i	���������&�5�����U&6�����a׷��w��9�\a���c��:�8�[*)���we���w�c�����m�1������3��6��P�wtZ���!�1��sVa����ope�w����ѿ����O`\>M�@NE��I��9G:ѷ�y����s����#*�o���n"�e+ް7��w�l��V�
b�w��촛����=���˸G�˗�$,j�x-����V`Ql|����ɡ�6�:[V���oF�n����e��3C���pp�?�/��|2�~���Gi��_)})����Ħ,w�f�cY�9�����n1��l;�-
ra˂<�`�+�p�kpŌ>*Q:Mu��	�T5�w�r�]9>��Ҫ�bx�ݚ�l�L�YG ��ϱ���j�c�MM�׊9��F�**m�i��gx��@�voe�{��P,�e<q�t�@�<��9DS�8^�y���y���+ř�2b�7�����Q~������&y[g2,�fe��E�1�uLUn ,8�
����Vn�m��|�_ο�@b+��@{#K��:�5����g���]��c�Cβo�-o�U�c���ҍ�Ւ��ֻ��P�g�����1�)M����q�/t�F��hU3����7��nc�e����/d	�o0O6{+'��W���*p�A�>�K�z�J,%Th0��貸|#�>IG�ޞ�L�i�R�BX���a��K�ٖx�T=e�����u�i�|�*�L�	��-�F!6KG�*�Ù�Ȫ�0�{y��@��X&�p���0��kto�$x#idVvO�&�'�S6S�U� ��S6�מW���!.�z�!P�9&mU�Q��Fmo��>ZFM���7��y�a:<��A��J璃2weϤ�Г-����������8��(�P(�9`�aaÏt�=�8��0��&���s�c>ʖl�DA"���Ķ�/����;_�	�)��
p���i��GiW��&TlC�m`L���;�����|Z�0��Nu�5Ga��P$������bH���*vf�N�=��=���/�H��y�5l�5pPK	cdVf�z��� \�ƌ/ю;�z��Z}3�$�g�!��OC\�k�ӗ&rI^��fˢ9�嚆ך������fk�q|ԕ.ύ��98��8�>ߏq.�w�%ǌ\9��-�?��KoZE����Fs[�.�U/�(��<y���R��EI1����۳ߜ�H�i�mȜ�n�Y$Zw�{}i&��Z�f���k��6��B8��1���<쾣��c�b��5��cO��$�
�x����f�d�U��Ʈ8�|�Aً]$_d����ǁ>���������ƹ�{{t��'ㄭ�0C �`��}������@�v�!�9J��+ß}�z���X�� 3�RN��h����cP��#�&��.a����<fY�����Za9��ϖ�!���TX��	�H��8hͱ��%�xm��U�I��E��ȫL�{�� �9��!=��Sߚ-��H+��(:�o��������m��(�:,hlv{�My�E��y[��R����Udg��H�?�26�j	�zc`�.�L�h�H���d�ƴx�cG=���fh�١�&����h��dl��Yd�b4�+�ܠt.����H�"*!��=�E�ͅߖ�Z��au�p�y���Xa7{�·D����:c�[�*��A� 
���aՕ�K�e�`_�i7����S��\}�r����Q�/�1�I�rVwP�-~[S�W4�����J�����W�r��v�
�/��s�hz����ɲd�\�>�ND�Ž��7&�1�}��C#72NU�Np���}��y��W�{�/�ΡbM���K����ǃ(f}{��~��Hx�J�78�����m��6Y�q��g~V�*�ݝu��g�~�>yKdT�:��U�.\W�� ѱ�H�  ,����j�{�)�<��?+M�%׫�����1]@x�g��>pņ���t�xD�2Y���!-�E�t6([�p�ɺ���pF&3Y�}0���L}�r&�vɡ�6�i�I�����B�Oe`ju_4*\�/�S<%癤do^�1�/�;���1{W.�wո��u��!�T�j�S=�
L���B�W��3��q�-Qi�dT}5���Ʊ7[.F������V.7��t V}�e>��᡾� %sH�Q#i��1B�'Ԃ��z/�|�@����q���(!��s��srRڭ1�����?N���(.��eײ�ӹ��|rr�=[�g���Z�/]IR�眾� ���O}e,���� 6�M��D?��{6ϖ�G�@K�>s�K�ɽ(|*]�CV��@(.7mU/�W"I�"f�+�qm3�G����ݝ��q�Б��jMU��+"�����'O� K�Zot��u�Ƒ#���hǧ���GIֲ"��62)Iz$
؋^Ӎj��6����zBĨ���2E�W�?��@�i�I�%y��)���V����aX�H�M@t�#0^�Mv���zˈv����<H���(9c�cQH SmB�Ќ��s�ɻ{96��j�CIn�� Ҥ���}��[���'�	 ~�*5���(�	i^���kM Y�6���1U�+�|:oyp!!+C;O~�)\��{ޝ�k
&(�l8C�x������x�ȱЅn�
0ȗ�R탽)���^y���X�]�s�Տ�U`g��F[��hx�H&zY��$�|K�<ٱauA�[�LC�Ҫ��������;�8�1!w<��[':f�� �}�wXB��	���w҇~v�%zp�Ђ��\�H��/��iEM�}g����h��~aݨl	�ϨMU���36��9)�3{�1
7�ؗW/^�k��6Y��=ʌ��&�b!8G�m�;�����"���x�Lߡ:[��\/M��ګI�sp�	�q������gx�};�%��䱀�9��]�v����B�C�������1���g�õV��+���!�2�f����i9���SȨ��>���&j���#4�L0��)"�s�\�3��
�[$L=k���#.�+![��?��֛���5�~Y�7�팈��p��ּl��zD��w��t`CɎ�IF6�2��~�Yo�Ur���:B���W��$��b�AΜj�P���Cr�B��Od�`�i.V;Z~1�gH>�r�!`�x�f�T�൶�%�6�#��a��v�&�|Vv7s�oȑ(N<�E`t�A�7"P�46�_&��e�'�+|x6+Kx4�o"�k\?����"�h�k�A�s�#�#�a�ޞrx>Ni	m#@%���r1ĪA������q�� B����/��-�U�XEȮ^,.H�0 :�!e�\X���=���_�@�$�����Y�q]�('u_�.��8�(h(!5�\1�i��k��w��<��ksK����o0�y01��������q �(�eL<`��\C�:0��f@��d��Pz|�;`��(V�|L�?��n��A ��iLG�\�~��	�i������p.#��J��&	�'&�|3[�7&��������ͪ��$4��r�sYm���`�\�
_�ġ�郎3�:��@	�[o�=���a� 	�./W�	y`]��ykhK�Ά: ����o��ط�W?�EI�g��}�*8Q��N�7�+��ל	ۿ<F�N��!]2�9a~�9���`���XO�Y���c�i�?Z��	v/���9ǜ)���z���Eg�+������"U���c��:k����͖�=h�P�h*Ę����	z�d)Qc���O2|���wm�TX���3`7���)�"1�>�˾�&�vq�+/r��+����tI�xؔ��\�����[.���~aԫ�M�����?���L�շ�n����� ��Z}���~�"��[��)j��P�:W���T��9� qB2�~.�b�l���)�����V\��x���J�{�"(g���~u� ��d�G�A�P��.����e���y%�Z�ܪ�ÙS�g���	��x�� G�v}�縝��nUWN&:��9������_�yw��/a`�T/�V۟ PC!�AOg�]�@R�8:1���>��{d<�|����{[���3�1��X�Y�̹l+u��I��r��K�|@~��5���{�3B[%�=�)럮�rB�S�:�xנBn�r�� 	��Ig�*�4h��w�����ZR|��y�[
��X�SRBlh�󜓐_���B��ņ�@�������T�������9��o�F�i5���[��c3[��=���9�*���)�4��C�evb9�����?
�R�7�W7�7�F��U�'�y��>G�$�2��u�pĄ7n�M:�|ڒ�\��9/���᳉���0ZT?+��#P�|�R@��>�/bۦ�)u9WU��>�D��s��t;�=`�M�������:?�3|å����F#�P���p���r�74��*�3]�.��O�Y���1~"�?��O�hs���6���S����^|���u+-bJ�zWfʯ��)"��}���.���Wq|�'�E����Sah���뗣f@��:��~�ߦ %\��;��^�&9D�@�����>�X�^9�j;LW���S�_}���:�����4q��&b써#k(-����pj)�ن[<�C�[�F�n�|t������8MO��L�kS3{���P��Z�$q{��U�۱���%`:�ŌΕ�����a �; ^^��w&��8z���z����!�0@~u��8� jdB5�4��\_�j�D���Dd;9��bP�^��5��C������$|�$����X��N1� /}�����"�=YY4�ʥF7F�H�x k(=M<v�Xy�
+�T� Dm�&�;0�>N�<A*�n4<@���0���\{�C9�ԟ����c�Jh��D�&V�W�u�p�h����IJ֐��T^���D�ؽ��m�I��r�0H<�$��hLs+\���!����Л��Q�aŇ�NŃ��f�ҵ�'>�/��f�@�ZF"= ���k֏����/bX��=�Y�e�Ӯ������xW�r�v�{��@�ڶ��O:^쉦�Q	1�5�9�zW$����]1�Ci�I'sX�ʆ_Ԑ��Ρ����8y����RYi������&B�@(�5�-t���^옻EHքz3'x�YʸkԤ�h� UR��DJ*W���9��i��) �+Eg�(^��R�p��Զ��o��Êt���|��"���F���C|fO�'������H1B�P1�t"~�A �R�fm�jk3�@ ɼM�Z�a��rp�I%�!�&4&vfW�xc�f�eg�z撖8�'�	4 �cQǡg��_~�v]�����?D�*���a|���j�i���~jʈO��)��Oc�O�>NGK}:�v���`��<�^Y���y/�@P��L��)��uz��b%	B
�9�/�8�[D�e�y��7`Ե�U���.�� oduO-�x�{[������ɟa�Ey�����B�Jy0�����5����!�	0��t�W�?�2T��y�\Eu�[�D�
�Cġ�3���H���H�� � H��QS��'�`��W{N�6���\@w{�|����4��;6��I���n�^�jfm�d7�������[r˹*Yғ# V,�,�3U�+�G���_�m�4I�wg���m���y���L���� yu��夼˙�V�n/�#`�.t�i��y�t|����*��TT_WVZ3%�y�p�m�� �飺Kj���W�] ��~V�1ZGk�W{?,H��h���?�?y�~��4�Ovڱ�词ǽ�j�.�{�_��A�E��B[��*�%��)u�A5&���^8�����]1Y8�/��f]�Q��%���KM&�V�������Ż3b�/z���1���a�v����d2�Qx�)�Z��N�( ���r���<@��P�XUV]���'[~եf�w�_�.j"߷1P��@���{��*���Z�SAxuU{���Ȅu^�=S���A�&��3�D�P8����4y(,ݔ��ޛ��{�Ko���gdq�����V<������+xo}���V~R��ԑ�O��ॊ,�$�������w��&���{N�X:���g{�@��:5R�{1}�r�ug���۔��PD�?�a�2]��Os_h.����	�㓔5�t��|�~1u!��Q3��Q`�wr,���?VE�(J������ە:�a������Y�r��f��R��}]��6l��>�����{�C
�
2�4i�����zy���ud����R:瘕��^��Y�z&��<'�*��3�|p�H��&[+�.v=�w��2��8 r�!u+�_xO/�J�e��&��vi��K�T����K��(�iI�՚{¸�}����� 19�"�Ú쭯�2M�6�z�eL�[�šT����Hm��:ܪ����O���@�I]��q�0^�[�2�=߰I�8�{D�;���p��!0-�u�=ɼ6#�*��ﾸA_�q�nz��3�a���,���2��K�>���IB��w4x�`(���8R�C��R�� -zQqF��U��Ȁ ���������$�΃m^;4F�(�ciW9:���-����8n3��9���x��G���vt��R�@	-ҥ���Z��Zg��b�`8y�v������+�����s���9��'Ѥ�Y�b��8�vm=9>'9��A�:萿�z0 �I�(`��~�V7㭙��J�u7��E/O�$e��5�eK�k�G�'�)�i��	  ��8*��}v�ZM���
��"�w
�k��(����P�W�Jt��9��`J����kG/�!V�[��l��j�<�"i�C\��)��Tm$גG�3�]��/b?bC����/�i�Fu��u�v�+D� w�h�M���Kb~��c2��F��I
1���u+c�L[���W��O�f���2X!���9�Q1�L�
*�~��[�f�c�1�|ެ����w��b+�x����펕xv�A�P
��`�+��H�8�@@�n,q!wu�Kꫬ�-D�2���@]�g�9�>���ɰ�H�0j�Ub��8�#�M�vp�$*$U�s�$�Ў�u��2F̩�8�)�8�*cп���?z�t����a�����V�k$�D�Hژ#ؘ��9�3:�/�dKڸ�+�5�cA�����\�$�ۓ�ax����w⻟���DU��7���U��Pܿ7��,�51�so��<1�	����}�V3T�����>dT�u���\Ij�w8 �œ6��}qm�.�0ߏH~;�_S$_�L,�^E�Mº��p�6�z�gG�R�"�e��a���c��7+�1�r&Vms$���s/���>�˺��ɫ��~���XRn�ZwS(�,�8?�u�(V����?��<�ޫ����X.�=&%g�ӭ_k��	G�h{�$a�3�ũ>�l��WEB����F�j��5���v)"�ѻ&V5�V�@�3�~,�҅LI~��:zi��+g�0�sAex�5^��k��웿�~���ƅ[�-#t����� O��9Պ��Y���7 �P`���F����L�q��	�)�F�ů���]�Y<��ح����Mb�XDC����F�	JW��y��
���-��N�O�C��b�&E�A��QQ�_��+�v���J������$�!]f�*Ǜ����<&N}�K6�����Z�"j9>�w��sl���'������-��}>d��:FlE�X&'=�nUT�#����",��a��������Ü��]�?�h^A!%�iD�ayK���1�l��1ȥ�S����V�%Ũ����w�mHO�oi�2���U@���(�M�H��z���$R�����q�m��_?En�=�ל�s&����v���l�6�C cw�����x�c]ٳ��=g�]	У��H@�.epE�z��Lye2��.�H��'�S�����AO��^:�SI�K0e1�z��!��''�;[����s�مο9�$��/���@Hq��n^�)Y;jJ��R�@B�^���E��!�T�?�K� -9��9���uN�#hZ�;t�Z]F��}�A�H@��4���}�-�X��W�C�\0<�q:�_����1�� ���w��uQv[�û	��x�����N�>>s%J��S��_�ρJ}M@�W�D�e��h$<�,3�h=;��x�B�nE�J��՟��l{?�",���r0�Z+S��ϥ���҂����3��q%���/�,T�1��w
ă�9+�`}��2�Uy"�j2�&�lJ ���s��`�ނűX�	�{]���l�%qG��M4�j�#,⬐z���Fun�?a۴�?
}9;ߚ�fV�|
O�e^�����`�(;�m$��ֽ��t(*�@!B�����+�p���yn1��q���8���(-�������zۆlZ����~�:�p��1Gg/�F�⎹��,��c�H���IY�s�8�Oe��n�`�3G�s��}�Ic�/:��+I+o[��dOf/#J��x$��\l�8UE��?w+�.&�~3��� g:"��8��W3�I�:h�ն/?����vz�e�}�/�T��	�>\�zն���3^xA^KU��
Z��e��~���p������!�0�\l��i�;a�Dk��@4<m&��eg/��\���q�@o�૛�i}�|�;ڌ�w` ~�{�?w�P�Ǚ����O������D�퇋���i��P�5g/���0�N����n�K�6�pl7��Y��;��yǼ�c{���{y������k� ������&k@�xP��҆3k�荒�[Nb�i'�b�
gia�GaP�8�j���H3PDT	���)�Y�E�['�ʝ�xȸ7���_!�Hf�	U_�G�:�@bkw������jnmL�4D� f�רk�-ޙ�4�'���7��{!��P�^=��oX��7;Ћ=��l}���_�}9 ���������b�����8���rUS��_x[Pk7�+�c} Ja��c�����n�j��/΍�l$5;Ĥ��/5=+Xn�]��r��A�!�Qg:]}Cg�=r-�l��	)%������a������ ֱ�>�Y}S�z�R�J�ƍqeb�<8>�e�7}+Ԍ�>��G��_Ҋ���ZpׯC��'��[\כ��r)�]����Cw٪r�@b�0�)�&�8�S�.��\����.`�	���*R��R�� 诔��[B�?����<e8���I�x<�N��:�4�����
S|� �'�XU|J��X��	"��w��K��ݣ��h5��?��`
�����On�Q�ظ���Y~{(|͵��=i��b\�i`�Cm����{�����܆tć���a�E�F�j�zG�_����mt��=u3�w���d�����G89<\zd�@�d��(WX�<]45}�A�W||��y|����ڒPi��e�H�{��s�b�,9dA���f#pZ4�H�9�;�:��Ԯ��%a/�tat�R��Y�E��$�9d�l�<f�� 1P�����<v�^9�(T�������\[�x��vb�U��+��a�<`ZwT	h�l�+�~��+��`�3m�,�W�k(Ge���#X4W�	~ ��N=�3͈��:�^��P|%	�bQT��s�wˇ}�ɾĢ=;�!<Lk,�]�Hf�P�S$F��0�Lk��)|Z2���;�;�I��#�+�h�t����t2�@�w�����5���Z�g�Yu�Ό��L�|lC%s��,��)߉J.���^;��s7H�OЫR.��m�W@��X�EpC�s/K�aH۷��K{�
�I���ѥF-i'R�v��e}�g����=��v$��;@2�}���q��G��s�m~�;��*�x���a,U��%������%��Dc�P���?�e�ڻ��|�Z��g-e(�a��$l?2��K�9*�;�Џ�Ǆ�;1�_T#ϱ�+�@�<� 4����	,c�yf#�<��T��J4j ����K���\d�#��S��P$G�B��7$�C��`4�P�&���v���0mƚ���Jpa�����8����,�
>����{|�v�?�'�T�c���q��)���R*7�]¸U�$,�h$J�y��������z�zٰN��_r8ezn~�����M�B�O�>��-��M3�'�G��f����z��A�-�q5�yuSi��U85_w��`{)&��\�@��Sn��R'H}e4I=��塬�k�:3���&c�_�'��s��y�+�003
��[�	�8)�^n:8�8u�k�F\\�����(��8;:��`�J��٩I笒�S7G:ŕF�NH,�mx�G�*�H����.SmVf��h'X�cM3�����,׷������7&ϲ���H�J��B;��bm>�ܳ��f'��QAUU ����.EG%�c�+#��[���&llFH�Fw���.�0���J��De;A��z��ދ������wQ/�̓b�%��oS# 'j�3�n�6iY�>���G&�:"�N�4e�X�+�FM���*MR<�L?oO.�=� >yA���ЙCr|"�z�6���tp!�*H⑼ˮ�,�Gc���]܃,ܬ��!*C�3EqA�q�W�uX����Y��/�P�ۘ�r#�m�4<�aw_+:
9�^��8�6�]]�z�����zQ�+MM�0�e��'�U��s�X��m�
y^�������wK@Ú�8"��#q�9�;�^���]<�_·̨ vLpk�Ii_��]�+A������C�Ѯ��v�˶`t��5O�cր�5 ?x��,�gw�_1qrK ?����@��4ЈHh��J�a�#?���%�_t��jin�i_tѨ��r���dB�,kj�ge5<�	�]�:��z�i k���I+�0�eW#����Ev1�_<V|�E���K��}?s�����iL�s�%*>|�!�8����_�|�Q&^ȭ�𿑗`��*�X����LN .�S�Fo�ܰx�S�V�������E�O��y�XZ���)�HG�g@�9R��T������/� ���O�>�a��Zf��z��c~��Ï׎�jG�X�s�g������>E�4@Ӊ�i��_�̯�#�=��Q�kf�fqE��8����]�h=��p𢫣-�>`���ڇ�v��욀���{;��R�,Y:���y�c�1i�޻&��eM����Y�S� �����F��-����G�m�^O�f���F˳=
�Z��`c0�-��P��sǡ1j8ʄ�2�d��s
�}rį��7.���ȴR�Ʈҿ�>�z:���~��7�˝�������YE�'��]�c���?\~�`h���|(%�~J�ޗ[�[���a�;`������G�Q��"�m�u�Vt �<��Y}w����2=	'�Ң��>D����f{��Z�(�Y�Ρ*M A.���� �6���?v��T���,�G�Q�y��F����W�혟�܎�wG�H7G��	�(a�������WԷ��>�sr���8�d�Ubs.���� L�A@M�`L>�zUSGc��&DU�e�"Shu�{�ʧ-~��gj,�z����k~���$���>[��Bȯ�f�׼�b� }�L��.�� ���i������Q$��TTr���,Q�&�j_�v�'�dJe�H����y`�B%W	�u�����Be1{�xH���<�/�tN7�� ���Z}��[���}����rn��8�Q9�$�r	ut:���d�M�Q�u�h��|<|���[<�>��^�B��\���sV�O��c�-c�֊�O��a�����qxʤ�6�J�w�/i���B����4f��g:-�Ƙ�k���s+�91 B�g��;#�"v[Es/��~�I���a.섰hm��B�h��a\(�|�&�\n���=��p�81�\�/��Sޏ�2n`:�ya[l';��>�+����zJ�纕'�s4=<'g�̔5�ϖ8�}��i�?TG�
�2�WJm�n���e�5����bc~ }PqY.�!bHEXʩs�3Y&O��$F�`EooPAX+}�l��+l���0U��T��R(�6�,>�.%5��W����4�Z���W��CN4�?_6{i&Eڋf"*T�qY
N�v_�ld�%�I�	�$f���d���\.OS}3z�#$�'y-�Yxj�&�"�2FX�ѩ���n�g���� !��k�B���Wt���>d���uO�ɟ
�>�Ľ�����N���.�2�����^-K�;�%�rێ�n���n�k��B�&��J��3GX�X5�n�Ϧ�����puN������n8��JT�2"V�:�	��چ����~�'�B>#�*�%�?����{|l�m�%�L��2��*�B��/U�a�<���'��圗��ʍ�8eM��)�Y<Ԃ�m������D��`�6�/��[�z�5q�W��F�k8��8�.��+ �N+ !�ڗ+��C�<& �W,u�#�`l��Ư��}o~�0������>Q�}Cƶ:_#����{d���*D-;"�I���ڨm��aF��ƾ|閔����_�U�+�wqCXw�K?r-KȾUK	0�PG�_NL����A=���o�0U����͇������W2ko_UN�㔻�@�����.��ۜ�����Z�z�e� m�����/����L�a���<d{f]�%�(u�\�z��f��Z��R�Y��+�%�.��'?R)q��?8WSI��E�c�{ʩ0�";S��f9N�<|C���@ؓɭ,A�B������͒ ''{�I�d������z<X���8�|�2����eJC�~a��0��r���hUu���皆�-$
��D�X��ne���|�<���L s���.3��;M�#��d���K�X�w����~@׹f�R�25�O�w�N����|l3є�x6��ϱ��)ϱtΰH������l{bP�pև N�E��'ݗ's��7�Y�2�C�p2c�%��ʈa�\ ]�p^�mK��UޒO�s]��v�Ǌc`�Y�4go���;<��8��f��rKбѵ$��v[�[8 :zH���۽f�%�H^�D<��jű���(<R�x�O�wB\�(zk62� �j���8t�5v�çUZ8�t+������L����&�l�a��N���ΤMy��:ђ�9b������X��9庵����p)�������Z�?��d'��$�H������巜`������榚�/�t8��ݕ�������$����~(3nft066\� � ���#G�'*?�W5�.��ěi���	]9b{�^���G�'!�ty#�U�?�[��`!U�8��i
&�J���LȂ��1Cu'W͗����d7#M�`ϋ'�M$4���s�%}��[.T,��<�z��KP"^`�V�m��_W�'�	ت�f�����
/5c��m�q@;�0�G�i.ݍl�&;BߞWq��|poc��6E����\3T�zp/��z��D�_X�+Xʟ��^C����\���`I?o��K�@��q����9�q��#��<�[6�Q9;ܙ��@�� Sl \��L�Ը�N_�A��5��;�"2j�F&�Z����QdD�m�;�˫1XA{�'�g�@`�j��el0�]L�}j��J��F�v���rXS��Β��?�Nh�qJx~=��4;���}��ׇ+���������%-̽�/��(Z����7��T�vP��Έ���	o��%mڤ��N�*�-q�����Ё�� ����@g;�d��M�# b/-����n(��X��4H��tih5��+l�6� �f����n�Ҷ��ƪKY�h����D��W�<�d�߬8@-2��uL��87�|��h~����i��H��+ ��ニk?��+�ӏ��6�U�o�o�ǅ[��,6$�,��`C70��G�[v$�����f�ˤ������GNl�g��k3q��U��q�vG��x�҈�t�o��Fe
�_N\�����Q����OEť<��VrM�N�A7tC�&�Q��f&d��}�\�Ŕ�z[���X9᧹Ns~\����D�gb^�5a��y��	��m�Nw{;�佼�
����+;�Ԩ��J�T�����Ə��YrP�o1�,<G˂�#�ʉ<����:�@�vi��C��ɵ7�o�<�(�%�,}�U[@޲7��X��fK1�9���.�؋*�L��#�Ր�E<P����Fz��;:�1rֱ�n�"��U� {ePGW�y13�	Q�ۮ��7 fNb��;�e�+��	v\�����Dr������rߴ�w�3����9��Ǩi13]��vdgl|p�{~�@r3p��|a?n�ch�:)s8}[�0�ז�I�oГ��d��mRh�[ HV<�A����'3����k*7Ta���N�S��ǮB�s�Aر�4a�����o��>�5��֗��ϧ����F'�j>Yh�<���:(���Z�|� ��g$��_�ssvhWSO��y�	:����3��K��^�?4ב`���%ؾ�ѩ�w,U����Vd�Ն*<�ݑ-գ��r�2�9�?���u�[k{̀�3��G�`��z},a�.1�]ȟ���(aBl�"��۟)A.��t����@�I�7��^����R����3�
8�7�����Qd���\ɉ�2����ﴐQ����Fka��A�iY�ȥ�]�fM�$�mZ��TV���J� ���C�[�v���9�NNJ*�<�R�����!��|�g cG���Y ��r�K9�쨉�_V},/&b�jπ���+<�'�3 �}g��N����ң'�U��1�*e�����u���avw2}�U�j.<"�x=�n*j1��_���q���9�#��Ҵ�!C���:���ٶ�[}�j��'�}a��İnm`�qc���a3���
Ԉ���5L%B�Gz�ú��l���,(XFh�E΃���L� �ӧ���T���ʜ���6�x=��Mr؈�4����H4�J8�6tp�Ǥ��J�$�&�/@0=5u�-�
:�����K��������{�p]`]�\���e�~@��.Μ�\�!+���pd��̟�%X����iB$=|x��<r��R����R�z�[�+g�'p_��'	��� 	N%�@�#�2e`�G�I����x��i{%���T�J���n�P��re�����:��Ou�F'Ux�u�8���j�G)q�7^'�}�����ݮ'T)��a�m>[��o,�$� y٠w� O�@A��%c���e�%��ŋ���7�Xg��d�t},��ߝ��a@]d��<0����n.VD G.�삼����ӮF��j`��C��Р���i3I���[�����C�.�馑<�Vu����Ңg�o��-�J�q�ߧ	r\��N�;�z�X�1����Kco��M����tx祌]1��{�1�Hr�<p����Ĵ�0�}K����kc�6v;��(��}��^�BpQW�H�i�F�2�ek���C$j��DA�X��ԊOtS�ࣧ;�$'I���N�ՑS�F}����r��`]��,�p�Ns�2�.g�J(W���k_��Y�νn>@m��"��,9Z�yf���kzÏ����A}�qi�]���7�D<u�JV�j[�9�^��s�����^�R;uqz�k&�?8�2�s�'�UZ8�:3�k����P��P��ub�8.��*a,��p��
�hB{)7������3��+��[߂ȂA�ej> ) �?Z����ad�!�8�9��&��Y�)f�?|*���=���̵ k
�sD3�@7к�իp񴑎k��Ǿ��/��3Xg;��n)��IK&�Jr,� !�y؞��4Dl*Q���Q��K�1���;ת���iM%q���xSﮰ�C?�-ڳ_���1wV��7�_���]�(�X��}��<p�%�sﵤ������!��g���XWT����^;døӴ�֗��!(��w/�"B
.$Vh�Q���{4"tc t*�7X����!OիBS*}���y��IHp� k�&K�SP�R��Kuݤ�y��dSHC��Yk��48#�ò�N���ؠ&M�Qh
�1��\����6��v̭�Żǥ��!�
-�J��Y�܃����~��� [�W`^��^�d���P;:����I��� 
O>�iB��C��N�bxQ����q�+�ԘT�C�J����vۏLj��f�A�$�8�ď�t��^ezcx�0S&���a| �J�7�u�tc�ٻ�����a��m�����~��=�D#�C8cQ�YM]���m����H�kS��Os�bC�C����L�gGҍ�֠�x"�T*����o��U�=��V֕���
�^�J����)|Ky4��Dƙ�H�KG�a��=v|�u9����t�,��Y@���Ś��J��%��)u��e٘�+���Z\x� �ӷ�M!6�)5���X�Ck|�@�������u�^�__��-eQ��#��
$�S`�3� ���ři�B=%(�*����z�`����z ��>9Q9�y�
�Ls6�֧���fD%<	��˒�r*�v׺��a�� �@v��Q�U���y���M �x_�4h�G:��ork��	��O��a����Y�M*��'O���
:*r(+�l����W�$Ү���KJ��,3��e� �R�u����v�M��F���#	��5���Z@���I$��`�	�w�`�"Ȟ�<�w�� �nt���Z���+&36Ɵ�']xY&�q�QN�Tu_���lg�U]W��o�q������ZF�ZD��IBP*�o� -��ک��K^{b̧`o��e���8��Cy9_�����6r[)��4IIYh���58����tDm��7�[�����.�K�B_�߹�:�iȔ3�'��px7��Z����
eq��	?2#��3��N�xd�c]WRi��rҶ&�Б���UX��dSZ���*m;�&��S�|<��e�`f���$������d!c�8�τ�R	(��O	�3��O��p�J�F|ˉˌ�~����$C����P54������xu4\V.K`�'-bq*�"�D�ussT�+��	�۞�X��#��1Ѳ���)b��q$V�_D�P�>?����/����u)�um��b�<6��&���]��c������4i�8RgC8�i�Õ%���`�V�x��u���?K<� �[��w�d��Oź� ��&䲐:8�}m�����o�|8�ə"X��}_��j�6���^�ۋ�>�R)����U#I�Yx��<0�sQ�Բ��cT�`���Q�ٕHv4�ǻ4s-6y�+��WEz��ƍ��[B��}��(k:�������Ά�|��I��M�]�A3���]�n���x6�֩*m�g�-݉t�+�������$a�x`}��O"������)���$İLc�MB��xc�����X����4�oLa��Ȗ��6I�GRm�����G8��x����j�a��j���&�ǦGh MQ��"�P#�
�&8
A���/�/�OC7't !�c+����a;ZХ����)4��>r��I(�޶vY��9�?�76�}ClO�*1��U	ȷ�8�����e��:������*̨MNLv�n�oU=UU8I>���nF?�q���L/��#[�J�D�Gf�52�-�?������U:�!\���ϡSnH������j��T����/j��I(S�6��B�瞈U27B�-��
�'��z�ĸ�pLuP�b��Ia��}F����
��l�e,D;�D;��17*V�C�m8c!��8��Ia�y������r�@-�D��n�px���0�f��������ǂߘ������>7xPqщ�ve�؏�o�����ؾ�1g�R kTo-69����_h�p�c��8���c4F���&^�/����`z�d*
�^�������~�-E<��y�]Ɏo��I!?L���2�{+���?˳�w�5Cr�\I%7�e���MV`��EB<��}�����d�X��i��W��9�׼R�Ĥ�	CP7�+������߈�M� �8��_}�$�;�'g���|v�H��L�3@���k��a�t������G����F�����^_��ty__컩OԤ��{d
�a	Cb��;��c�3��a�͡�	ȍH�
��c�.��F��nZ�b����^��CY�DK�?�p	(��&���}�G���{gjd4�H���(�qp���6�]b'K�ޚ猗�s7E��*��V��d!�;#k��͹xE�JJ8��x�F4+!��Օ���~�c�d	5�(�yCçȚ}~��Q�Μ�y�)ː3�"��Ҋ��L6�%Ē�yE;�� ;'bF������V�Q$ՕQ����O����^)�9zPB9�uL����C��G�F!�ł;.���	�ѝ{��]�Ԡ�����r��A��HƖ��v��ZK  n��p8�C:�ܚ����/��/\2��q�#?ib�c�	H�뭞�X�0�zG��n%Z��Q�eO(���1��{�=�D�:Նb��f�荤�\*p�w���K���I����E��}�Hل�DѨ����<xA�y+�w�SY�F��s~��F �C��jO �j}���D�؍��ZԵr�`R���T.Qr�8��Fx�^o3#Mw��<"�̓�Oq1�Z�ۛ }�*1E�A�,�-���`ƿ�ٶ=7V}X6!�2�y��M�����t*��}��	��CC$�0��X-~����Wn}��p��C�'�����MJmɉsmY�ƥ ��6��������[/ڝ���Y��2"�o�X��s�%+˗ %�Φ�mG��`ؾz��c�;P�<���>��/s����4�����62@�n��t�a�ׅ'��/�=+z���>��?��J�|D�����$��H�t��i
�u�a&��-o�F�㒗��������yZ��Yc`��o�bFCu,`9iݯ� �m��f�����AQ��,f�n���Ԁ�?��m#��λܫ�W�=��D:��xp�y�ׯ튜k�PдL�8:�� ���i���)*��0U:�'3,�7�b���hد�#]2\R7��/� ��U��Ƚ�[� �=�l�u(V<=��!'�΢�/|�-J�M���jpI�LY ���%���P�Y�V�����\�#dR���(>�Q����;�Y<��. �)/���O��{1�jJn�ƹ���k���C�j�|����2h?�=~���q|R�v�%��+�<^d�`؏�lHF,�V]� چ���Ƈ���&�|��o2���ҿS�.M�=��C̜6S3R#�) xl��*[���L�+G���S>S��9Z�H��������Ru���7�X�gz�.9��(68rN���Iz=�6?�?��}���S?��66�_���	A馢I�N����4Q��2ZɅ#�<@�1�����A�ޫ���K��Nd�e���؃�h�@�e;eǇ��N;f�t��KZ�{��?H˸Tx+y;eila����w�u��Y���Q����\>�����+
�.�'����ܠ4xrMA37}�V
)�<��ﵬ��N��9��ugw'�eV�|2T�´P��+g
@�]	�[��d�ĩ�ч+�u�/�[��IG�LrL�qf�v�W�b�j�ڧ/��^P��t��z���@�~��k�yFB�K�x�e�u:3�LC�i�J�3~_��*����%h�����a�)�Hrzt�dM�=l?�*$�v��\�-�x$
�"�mЫ98�1E�)��Z��Bb{�4Vm^�#5��@(zbk�X���Z�kz�0�K\]/2��.4���:���]�ɂ���)W�o-@>#�TP<�\����Nae�X�$�	��̤O��ͯ�u��z��h�)�*}K�!	B��z��Ě�.���@��Ϟ%��8ޟ�K��?������T��i��o�K�vہ���H�i&�qL�")S�/��R~�Kp�'a3����}*��P�5�[j���]ٞ��}w�
����S\;9%PG�s᱉TcR%��t�u�|g��a_����?!+I�q	Ghf�Ų4fv~�?L2��i2�3�%ފ�wZrgs2_+����Q���DY��Ȏ��Q�u��^i�7w�^	#���a�0��Ԣu��g��K?mK�_�
(2�1���l:6�v�~M��&�m��@��j���"[*T�Xz�P��!��RV�6lw�ͧ���2�Uf�f�>��k)Sl��i�.��:�/��ԝ�R���ѭg!��oE'f��E�9Ng
B�ÖP���+��#\Cy��P~���#TN��m��H�]�������'5�$��x�C-�X�Η��T�W���V �5A&k��ٸv �k�j5��T���4K|H�i�� �`}����&���o<c�}{��w��*W�u5����r1�e�-��`�w%��XL����#��0�C| Ą�(C,4Al�0��˺�(&����_��k�3k!z��)�ߜ/0�~�7+|����ڤ1Y|ֈ�A��~՟5��qC��m�~??lN�S���7"-�#�lL�A��v�rrq���3��,5Ē�M�u��9�<$�!����^�z���d��Ȟ3Js��N�f㿦�UV�c>%��A����U�RY,q�'�5;ρ�m�#�o5��Q)��$��v�!=O<��k�@�� �S1�u�~���[��q���߄7e��WH�M�
$}qÌJ�ư���iq4j�!�>�x��̠�E%�MM ���K4�2�!@�.?$ �N��VG#��D�U��y{/��E]�
���Y'�[m����#�p6Na�Y�D��7�l,=��/qMɮ����n4��X҅4�}���H�c+=�rI�ӵ�]7-��[��5�,!�f��a<��$m+{xy+�����Z1l�m�"�H�W�nGp8���|� 4���z���-��/�U�x�J��l�����j����Ħ_��g�}i��2���W���d2�E�����#w�s��\79�k�Hai��C^U�H��#�+�Ă彠��=�v)�`y�LK+¨Ѐl*�Z=�c�b��� �f��¶o�JB6�{|��x������zT������H�An��e�O�*�O�R�g�i��X�܍f�dҍX�Y�n���M� �N�N�M؛%�SL���guȃo���v��/��Vb�`*:���g��z�nn��'��z��:�hgn�T]���"c�z��+�KJop�k+�a�&�Nť5����A�<�w^n�|ʢ�17h�3cZ Z%�.5�=m��3#֎]��p]���<�Ó�f�����L��D��sZ�ָ�a�����N,��7�2>v������9$E�7%�\�س���n�`���бOLY���zT�z��a13}6L�܇Z�aۥ�Eʆ	.��I �|R���аrQj��s�o��Ę=���d1Y]2�ƍ��4 �	�;
�&me$T�X�n!����/�5��AM��`fA��z2���Sw��Ҧ��8;���4:�9=!zwס<����'cc(�]	�kЬ�73�k0ڤ��
��;�ﶀ_/�)'��8r��갧�˷=�A�������Q`r
�����`Ҷ�E�d3#���E��B��8����]��n��@�^8�)��s�t�n�|8�8�ۛ���������dy����dW>��a��݌V>��.9�A��t�� �i�խ���ˆ*��|��x�����5io���{���'��vYJW�c����6ؿ���;�v�-(ʸ)ro��U�爦���2�*�IÜt�ob������/C���ir������܈k����F����1Smߴ��c����ɥls��-=hDZZ�ybY驊\��.��,�L_ Zp�������"?1�$u��(>��/m���-��6�yQB��v8�WF�o�l�8�5���4m5����J�=�C<X��T�u�,�� ���5b���N�2Z�*z�,X��z�S��"M���XY�9g���8Bp���!m��IK��Id@1�?��dI{麽��[��9���.��/:�-Բ���0��5��1ŝʵ�,i*G���a_c닓i�H�\n¹���W5Qt�"�.t����W�����T��k��ܩ�g驎ds�Ԣj���$;�c���B_��Z������mԷ�7cD]K�q@��9�0k�'������l$�k�|�򷒇�3�!��B�W�ۨ��U��^o�G�������d�:{׉��Xt�}r����m��~`4t$w�B����g�$A�O�u6��Rkd�q)���L~@�uoJK��l��F���R��i�o�G�^���	��Nr�{u�T̥`B��x�VI�3��!���|��/Qcʏ`X�,w�����ΛCj�X��6��AA���+A�=Rij�>�� �O�"�%M��5κ�����l&���LJg�Y�Nu�_����*�x�P1"����3��D�U�V��Sa���x4��s�ʬ-P����1x�7H�i{����}#��{��1"��v5�,XUO�!OƱt2.k�����N����Lg��:~�Q4�K�g���f�7�,! DT*�cэK���ўރo����i����W��'ģ�]�G�0�Vb� ��k�^1a2�7R�}����Í�C����7��7ݟz.֨M%(���d�N5���9�{֋N��t
AbB�?��1.T�v�3l��AU��XA����kӲ��%�'�a-p�=�� �~�� ��*��to�S��5�G�0@pV��0��?^�<��������,��I�Z��6(�� )���Z�YI(9�9��)jlL�e&���	*�u	��ͣ�8�`�t��'�������ۑ�<'�U�V�f\<�LY�T�p�5Em�w��-S�UXܖ*�q�cs��>n�huo��l�+@��LvIeF�ʴr��CL{��?�cV���d�3��״�'��Z���(rg��D@�*xVa/F����W�xޕ�T�MT�	��}�+W�I�^����c�~r����h�ڽ2��1��X����8L��L�q	�_Jl�)7r�k�[��|b�͑��z�=7��������2�,�x9�|�{�u���O�� X� Ζ�B)������db!�Mcd1uLW�?_'u����ls��k�����6�Ulw��o1�p��RO7&�a}?($�����m+��|`$�/���B�G��bfN0#�y��r���E�jY¨;�yc��TW$���e�@�z*riW`X=S�R_f�����0v��UVȰ�i(��5��aӬ隱�!ꃿ;��skm�Δ[eP34\3ZHĮ6>�@�?!K����k\8�Oo�W�r]	B�=�5�
ɶi��kgW�j�d}=�~�����8��m�'3�l�>��!Aq��S���+�>��⁅����)�+gu��(NrDX0�(�Xyȟ������X��{�l���cĎ��H��G0z!����O�h��*<:O|lg�������@�^쵔�� �B�Lj�����gfZ�1"��ƽ�\�����b%���h��Q[[���ۊ�x����H����a�[���t�.�^�]��]�y��F:��(��V�cg����qc�N�d9���/�<l��P�Z3���ۿ����#C�ߩ�R�#�MaZ@�0}����@�$u�e5K�D��}�%A^tו�3r����D���F��
�r��Md&Y�r��P�=��;^�ӝ}M��aoΠ�(���i�<@���(;P����=�F��~-�fh*n�r�2j�BO;~���-��_il�_H�,|�[+?�$�Δ"#D����� �7�<���y84�[w�d�1�
T�����y�'�φ+��u"A�SXh�����<G��B���>X���QA�jZ-e��&�YU9Pk_�53��zK�D=��U��֛NǦ�r4o���u�Dg��>7	�` �y.Ӽb�����'��

p��c�Ȟm�ͤ�Ѱ0�]�g�B �S!�
�Ӝ֢A=���dp��iN#, ���ND��x��H���<�&t��h�~a[��3تpj�:�K_�eOϸ���=�.�Vm%>P����w�K��~��}�D�ǜ��k��_�1�~��L%��*�h�/@�WM*��c�32O�����9b�s��	��Q<��&W<P���p�Bv�����\2R�Z�s���ӌ ����Das�Y�
��Uj˛��$P"�������@C�b��Q���Ԉ������{�[8�d�n�,/*����1�-�Z:�Ѯ�>J]���� �4"�<��d*Ҷ���i�O��.C�D]tOG�.Yq39)H}>�Tڨ��#�֞2U����N���Q�4HA_������O�Ս̜x��[�Ůsl���STl9� �Ph�	$�dΜ�F]��ɫz�\��X~�*6�(]��ѓutF����[�e�-Õ#޷��}�&�\7)��gꚬB�֕�ay680מ߆XE�?�%ID��YN�;Jgo��EY��+!�{2P%��n�9xp�"Q�6��\�(XS�/Rx�.����m[���@
�x0��rU���W]��~����J�a�'U�O��5�3;��,C���a��a��r�yټ����&��q����pb��ˇ=�	Ѽ��S֌��V�?)��DLm\�ǋL�Pk��a(Џ�UC�!\�IK�n �۲����.vL��Vf늩ʭ���׀����nmA.�0DO[�)�>F���Vm��U�u�>Ѩ7�9ʕ'"�B����B ڪQ��4F\���V�Z.��#��фL�c-A��mZ��F`�� �Ԉ�r8{MO�@R�i�O{�^8t;s�0	Ce����&���L�$ˎ\�Y��y�D<�ё��d���8�㒳��i��+ O�T�'�UePH}Ѵ�46�Bg9^����Q�-,e��o��l>6����V!mU/:f��δ��$*�
�)���"v"G(�X�DEj�wl*2t��#|0_��o_E�y��q���Al�ZԠ�]�s��\��wŰGH<�^̥�鵱�b*ڗ�8�!X�
P⑱��K0�����������������;`\R�f�� #���[���Q��DfMq�� �^��N��{/r�տ���'_�'(� � ��*��I�lEqT�����kSb�O�0 U$2+���x�X5��iм3�eY�&s?�~����D�WJ*�S1�^,�����{�^�*{���⺢\:���W����p	Ec�E��{�b9��j�5F�?����u����?��B�ߤo�^��98�B����Rt�mT���6�}(܇�Ѽo�zRHxk6��q1I�Nvn�Co�K�x��v�՗���
g��xi��z�!�JO�-��!vM���)�Ola8�V�R���֣�ͬ�=�w��Y�e��Fw�D�MBe�7  �҉�}Ƴ��0y�j�?x�;Q�f�.c3�,)�X���Qo�
O\���:	P�0�]Y7
`��@jtp��!��I_a.�:�ٌ�|=bC���q�������/��r�B��_��!�|dr�׋v��d�_9Y��X-ê�W������j��s?B�o@r�[T<�`��PW|Gk͓�˜f����?�ǁ��$"����L��W׏��M��:��e��מx���oz�49O���;���}��T��tO�; g� uY	^��F���F�	 ��*%���A��~އNXy�m4�R�wΥ����i��]��g�f �H�v�#�P�Z+>�"�͆�N���o�U)#�xU6O������^T���9���c�/`&�MR��4}�ư�ˣ���(6Ryu��L$$�L���5aXfQZ&�i�<�l^��K}YMM}�
@�7^9��XT|���d~b̤��X)^��Ce�_�&e�U���*�  �� 4I���5�nRQ�����R�p��cA0�K?7�HS�����J��p��Aǯ*Vb�-��A�gx8�i��1�����Y�_C���O��"�w��a��@����=o�`��E�uvF"�Zh3(%{~�A�������RK�����+��XY��9eyk۹�Ϋ�o!�R��æuk[���p�2l�R�����)�BBr�.�K��2���M�`ⷔ�*7�$�|�Ptvc���fFe�q��p�(�������4d9�>�hR��+���B�CC�@c�R��J<U���*x4�=o��z��wȋ�ʊ�b���	Hh��-��>���zF�G���������!w�	%˻/cIV^���n|�V�v�f͞c1暺?�E;y�ǂe�-sL��=�LDw'fj�8w��]!����Ĺ.>LC�g!�l���sJ���l���4�O�lh�����IܚB�z�qA���X�wr�!�^�R
ʀ�һ�Ϫ����
�rD�K��O��Jy t�fq� R�<h\�= I��pcUۘ�5��,`���tɸ �¸=iz���\E�bs��Mҷ~g)y�l�_�wyx����+A&>/���=��z�?0H] :��/o2��2�RK(�`k�[�[��r�K�n!��6d���+_�xM����C��K .��{�2��η	��Ż�XQI��$NM'���6CxJ�)[�~�Z&��j�`$����yJ�eSzО�1C��	9�2Υ�U,vG��!�T:�[$t?��� e��MC�
�}"
��8Ԯ�$.�u�f3��V���<N�y0`�ج����'�|�~T��M�U��ݲ���1;��[:��ISљH�-C�y�����%���ˇ��i%��Qx��e$����^`s�
�^�uO����eEl3M-��нN~���b�Ro�8a]�����t���`4�I��#:�
�3�M_� $��`;��4WH�����p ���ztG���>��,Зu���d����G5T��;n^��9��7�G��Ox�\�)�"� +�F�P��&u���P�O�ݙm߻�2�J��Blm�<��ǯ�ly��B���N�!��L�N�W���9u�t~Yz�R8�:��\0H[H��u�f���ï�C--LRO	��4³,�Ns���d�j錋��6o�R��*+�p��VG�up�CEebs%w>(�TMDX$����o��7�D�_6S��:���{t��$w����Μ�'MC��,o��;�ptF��.$��&;S`;���Ը*&� _<�	nu�&v;r��,�̸�wa��nm,��<�o��{�����~�@P�?>GWߑ"6�ÌlG��7=�#��@� �d�J�%�wUJ�Y �X�hWpքG�Ӯi��1�20�N؈5�{o`��O�R�=����m'�������M�O�NLԲ�$��Pm0���I9Ջ�14d����+�2��R���)i?��\X2?L�IedOww��<�8���pn�n�X���$"��:a��x�`�-��oW7U�Ǆo�kp��0s�����H��{(��З7���`.>�\�o���n@�Z��OqŜu��j��s
�s�"54۶;y�(����=.��E85?g��0;5o��l�e��y9��1�c��)���"עA��OgwKc_�J%���4ʹ�{��G���	Ŝ6�G:X�an�U���_�`	��<Ny(_�e	�:w���C"գa���p򔽞�	4�C��y�]e|#��\�V=��Pv�,큌��{@}n���3As�\5����%Tf;'X�RY��{��5>N���g4�	|���21}r�x�Y|rr��ϲ7m�����Uzt��y�gxqC�k@S��.��s���<��W�6>�n��2Yg��r�ʴx_K��;�mWd�7dl�4?�،��O����!Z��M"��%8�Nw	�ȠO�\�1��J]n5a�Tc]l�D�8�D��bzlɒ��(Q~�lT��	et��]6�y�/P�"NwGV��Be	G&eTK������s���{�2>Spr���_���(!쓑ϵ*��ۖ���H����g�B�+5T��$�U:���C��?��,b)��{��4y�Sb��IT����	�U���C��n*��]�o�G����nV�ۺ��[����mv^���ȭy�dV�L}��:��e����b��jЁ��S+��{}nB Ë���	������q<S��V�Z�LdԌ���?^"��|;�Cj��2�6�CP���k��C�`|]�u�͝8T�~l�e	�(��2��,RQl�ɜ�"�`�Ѵ]`�/L%2v�{��J��"4X���J����螏��.�@G��Q{u������+H�H~Ir.�t���4�!��=*CֹG��o{��iH��wST�I�q���}'�ڬk��x��"_��v�)�rO�~�sP�+���ۊ�W���J��ff��[�q����hk��Y��OذT~'�4����o��A�uo$�"��(�+Y=�tZS�!�>ه�x#~>]���OP�+��Y3�-�eN7�V�x�2旋��Sl��b9��Їr�|v��<ڈ�r�3j`����غVBFq��3��*Ѳ�i�af���P�<}�� ����ݾ��ǃͫ�
��tQy�WA����.8���F�����p�9!,T����|�	���z%'A-S�l����ra`���F���#��sZ3C7b�+�ؓ�h-��=w�8���Y�Wa�1�#��1����4�蘥���WK���q������zB*�XÓ��P5fj�Colh9�7|��z�W��ɇ���*�3hu��u2ʣ`���~o�j��9�b�TlG��/f��α�"I:(����]ȷ���LD�N�W�KH`�a��a~ʮ&��'��g4�K���/F��Cr�~���հ]�o�7�7]�~�>��r/Q�+S��Fk*&<ʣ��RÒ��r�jI�CZ�G�7��=���" m��Мt� <�k`��DCX�me\�������bF����a�<�;�GI�ų���2En	��!���`�5	Į����p&�R�T�n�O\�t�>T�P%,���.�z,���	���Y�|�0^JES~P�� !�����|�V��H�*����V���D�I�3_��ӕ���O���[��-���I�~�a)��kkk1�CbFQ���3��O�q�0�*�*���k՗6�ۭ7���&�Ev�g�WˬFȨ�0n.��I/y)�遥�q/��wmg�oU��UӾ�Mu���ou��N�(�������K��6	]�5I_�_����v?N���H�)ԮEq�p�I�V/+iP߼]Ay��;Ї����9��jN�E�KO�&�̚X��c�l*%q�׺,t��:��uP�	��2h�J��$� �-�%�ݒ��e�,��-������{ջ~�o��g'��tGN7�֩/���Ѹ�U����H��o���a/�v�܆���5������˪���0'*�[�(�&��5�Zh]���Ʊ�k��m_�ȃvJ	����Y��]�=;�n�q�+v,�Mɡ}%��x����$B��T$^'��N�w:�����F�����W4Yэ��A����Д���B7�vh�����Za��s�*��t�}�š�W����pcw�� �'紬��O��\�sU�i��D�x�l(��w�}~�ٻ��Ε�ӨÂ�U�1ʐ���=�5�#��+�u�pE�5Yw?Q�����*��(͆�"Q��[�h�����N��h�l�F����٧"��߭��a���B��sG�l����]��! #�w���a(H�6�6��2l�8�6:�&��~V!�Uz!ɲ�o������̛�d�ďI;9.�w֩�3��f�r^'��z��p��:���`���='��O��7�h��WQ^� i)R�}f��/c�(V;�ɒ�jh�D�!$�_�:�"x����)4�><�Y���_��+fwõ��-��|G��)Nz���1�=��[*�����:�������^ �$y	�o���y7��vh�h��`�k`R���.(ˇEft�ʫ���o#�xŴR!����]xLTF"�L���?bX|����OW8P:M�Lm�ϼ� ��#1uW윍���iw���Ӻ�4Y���&��Q��@�������{o�i^�}�gg2��
���B������*�h��UH�	#�IwS2��l�M���7�D���N�,�,���^��x9Y�"���W��j\��֩���ޫ�z4vXAL���7~�O�ӓA0T�����C\�Uݜ���;S*����>Ë��9���Ⱦ���@#�񀬚�����Vm����E��kI����e%����\{�j�y3Ѧ(��	P2�W�F�B��j�����'�x�1z���{-1�0�e �vK�4��c{��OIt�3%jv<����ɼ���A������h��sW��s�>�*0+���kwFr�<��U$_�Cb�%4ˡK�x����9��;2��s�D�#g>[�v1y�^[sԱ%�8�9��s?$"�R�1V����^�r�L�R�a�%���5�\Wۇ�ղ����\"c�Μ<J	�l�d��2o��P�)� ����g��$�B���V�T���R�s��� B�ѽ\g⢺>����E?���K�a�Bu�L�4��$�A�o�:�Z?�x���T-����w*��^������J�\���ǌ!>ħ�X���V�d��3�c�@Y�%${7� ��z�ʊ�3�of��T��D}H�.r��&(ĭ������Ѫ����ӯo�W���rl�L+�:�g	S��)��to��D�\͸��x�Z:��$���Uצ�RQ�s���b���t�,j*⎽��iZ�	��oB��N2��/��o�C��Q��H����9.�^b\7��P�l�v�^��դ���)�N������wm~B4���ѵ�����i4ɛ65�Zc��s�C�~�0	�i���l�(�i	�@�/ �����m�`��y��,��;{d�L��h����8��Ľ�^+(v��#��@�����SQ'��K� 2��ͣ΍�w\n�b�Sj_W�&�}��oy�@��8�C�
�+-N��k��x|҃�^^��mnB��c��ݹ�t�����b�nAgb/rF�YO}oxIw>`�d�TL�������</�K����y�<P둽X�zB�K9�Rvd����0~
s�ڗ���a��8ߖ����f�%�Oҍ� Lcg���M�G}ٺNh�,�{�����l���F��&S��!ً�J�<�d�{�����fxw��j��Mo�bg^-�Ϸ����VOs"��np耾�jf�/ �7*���b�3���k�.n�������-冿ِ�Ӯ�ϕ�FQ	�w�\3�*�,1`�<[@�����;ѱW���@�0�CYW��bh
H�OG��5��wx1F���$
l����;���_�3ILy��O ����T�(��Ӣ�s�ޥ}�������1L(��}�]�ԝ=�mwVe_���hi�*z��S�G�:N���6v��d6:
�rt�39	�~�tV�ܹ����b�e�T��QI�Ƴ�?:��] �Q��W�!�:��K�p$����8�"�b��	�@v�N�2� ��W�b�s��e�����u�;�O��l�I�W�$�i��%b�v�*�wU;�* @E�I�NE�@�mK�̆_���?�WW?o�.����#���"�������^��W�բ�b[�euƘ��-鐚Qł[�A�箸:&��*tDT��*��3��'�er��]�c�US���v4$�K�׵�~��:���p��ma�L:Jf��V�����X���)rTwro��o��C����2���� a>x���"�~TM�����dN�b��S?�A=��?�޾Ǘ�U�Ч�ZY*A��5�`���ua8㛐y�+�F�����([ںX�QjQ)���C�]��m���]�fPQ�#�R�ܨ,Y�L8�ՌC����������2�:/��[P�Ĝ<��]ֵ�r"(�}	 ����DMY�\|���}<�r���kN��{�[��j�=��q�|g� �4��>��E�~�y�N�����_"}�Eh��F�8n��P U�t����_�bj*����QQ��@�`ܜ�9����}�E�i*�c�&2���c�"%6!��k'�R�+����t6TMQ�/$(��8�K-P�(o�ŲW������'R���*k�OM�fGN��Y�1�6w4�ɨ�,��{d$���δY%t!I�l?E�OEZ�jK#TJ15*�$mN0\[���Mr7U<�2�|!8�3;WU��dh4F��܎���3��x��K�f�~A��CGa�Mnl��9�`yus��[��bY�UZuuyB��D�?7��0ڐ.yR�?�;K;��CȏdN�s��dG�����6�➖^d�I�_�޲�$:���EbΔ���
�~��Ld<�`��V����#����t�/�È�F�o4"���+��X��pix�{���_?��m^�c�d�������W�*�\�H���Ʈ������!�X/�qN�L�]����I�����e߶a"91�g5 ����簧|zN�'�q/t�b�j"����SL��r�{�X���Ak��/Ee4;�Ht��
�k<�c�u<��#Hyl�}��:�<'�h��pvxժ��s$��������
NB��t�m���b6��x���Uȣ��������/j��6�� ��B�ϸŷ3��%����A���3A�����-�����-2�$�n{���U�P
]]�CG�_T���d��8�]��`��h������;g�g�T$t)�x�b��.q�nѺ����s���L���F�5θ��a��G�=?u
>��m���YG��]���<{��k����n�{�ɏE��=R������P��t������/��W��aɔ���@�K_︰?��V�����6���W�1ڵ�}�C���p�u¸o�h�Ep,���OR��$�Jv�� �݈�O��&f���<,( *vկz�l��9\Z
�|� o�O<t)�%�J�U%�xɺ��;�i��d�Ӓ����r?�Xx���O*�v��`|N���W�zã'�Tqy�(��k�tHN�y%�au|v8�Eŵ�1D�H2�Hm�eJG
��P���}7�ˣN�ޛ��_K��RN"�͂�{����(�SyV	^��qH[�{������.[n�Vs�p���9OOח�lF���b��*ZV�td5��{���çr�+���Z��W �T��8�w4.��+*����d��b�8F���>T��@�v���'*�n����8@6$�	�W���U�:�ݮ�V�������m+���ү������a��u�4�t6&4H�u�4��9���Mݬ��w��Z/���QJ��Ԩq#SY0��8Z��v��?�6]�N���� N�Z�v��
 Դ�y'm�Ȍ��jːH��q���ˬ�\ ���Q;,S/���:��(��F��fFˮ"��<�]�"���;�따R������w�<Y(�M�1���3�
�Eyq��&?��*X^&"Y$@&��e���Z�r>��2+�v�<�F�l�ūb? 3�]�	�Z����]��pX{���ӷsІ䧱�o��ݰx5����$e?�7~�u��n���[	`+>�v�_d��m����19y�8�uF��B��������_�9a�x�_�s�D�{�`X8s�A�`E�5$]�C��|C�Z�#Fn�dX恘i�x�pU�e��.��oč��~����G!@P�3�Jjт�t��߀~��Q�"A�|�^R���K���+N5���7"T6{����r��Ч&e/�����G@�Q4��b*g%�:jr�Px�꭮x�(�dD������w1?.������;��1|���~!E�x
2�?��d�2�}�c��R�+�!����}�����Y�/,$B��I-$�d���Yf�&�83��͎��<��&O��J�/���hq��3��V���HIM��MkK4���ѻGY��$?��"i�*��$hA��#��.~��7J�F@�y�s���7�o�����w��������ΒlvJ�*����P-�p9l��+�Bw�uh�%������������|�>�y��]�AX��翛xI��DT��G�\����%�ە���'&d�s����~׎[�-�ф���F� ���C��C$�~�oi�����*���,&z]#?i>�&�kn<�ç��\4�l�����v
����	G�e�t�e6�� �dv&�?^�^>�&'�0�Q����)��O<Tv�5�6ȶ���Cc�`t
>��t(ͪ��>��h��\�{�Y��������$���A��� �Ka�TP�xӅ��0=���Da���p w���^q<�%�#���=�����W�yQo��4pz��gs����,kF���O�ˣ����ϳ\@nJK�g��LG��Sg��VL}��J�"����+K�dx!M>ef	�1�&��#Q��m���pՔ��3}r�)M���ɞ�/F4���չ�s�'���zJ2��<W��#V��{y#t��S��8p�Ǭg���� ��#�^�����\K�������Rb��j|�A���}KP�9hv%�2���J�{�y��q&}%�\��A���v��|�p��-姿?�%ƫ����O�8�����]�Mz��)+��IxT��l�\�v���9i\�	�`֊hv��.e�l^��!!dF7�H}�W��>��������=mQf���Q����8��-����/�;����F�9��֮ ��T�?4�����M���C����;��*��\Z݈��ki_���*�M��9����-���5ڐl��eukQ(B0��)�䎦���f���e[�:�
�z`�����f�[�����)#E>��b���b�	������ӿ.�;�MD �kz��Q0B%�f�H��3l~b0�����r$蒺�O�t��]+��i��|H+U!�d�������*d��0Q��@�p���op�����ک����	[�@��$j$B�_�Ҳ���kٳ�)ֹ�As�}1AL�s�T�{��v�!����z����rm^�=9����FV�,nW�lإ����1�;e$x@�
J���XW`�xM�M�Vp`˕�xO<�r����;���ҳ�p��gV��'!{4-�/������/��\h�b��g�"�u����d���'	��?+_i�ښP��¨�"�ߌ6-��Z����MD�쎹5��LCH$��<��	i4����(>V�	�6k
w���)�ۃ�Ťf�@�� �O7b��l�m�rz�دa���#�<[�7�a8)�7�|�\��~������U%�� [
=��oD0bH�<�*�D�>����� ��FӔ(�Ջ�
u��h�t"*V�k�q0*�'���b� �KBb��:�q϶3Oht8?⑰�d��<�� �� �?�D3uC���%4Ӕhʡ�Y��A�U�� �iqk��e��1-.=z��?Vħ�<]��z?߫$���TM��A���hc/��eȈS�,�^wl�E͊�Fs�+�@��I�@ZI�����ID��&'ʿ���C�������M)�͉Q�k����yA�D6
�qE��Kg�a��.C�����/��Wĺk�%�T,=��I�9����םj�����'�r�<�㼀 �b�߳PHs����%�>�!C��q4ot�K�����9]���6#.Xu�+#��3`Xd�Դ���5A÷ZT�(�x��)Y+F�ϷK�I��n��SN�Q����祔��ޢ%~��'�oF�EF P]����^�KC�����y��cO��5�e1E��Eԧ|�Z��ܠ�C{�u������8�xO/�858#�i��ٛݟ��)^�X���8
��_�-x�-X�� �dꭒ� -oR}=�J�l�/g-����y�^�48�8^6��j��\p��ɀ{u@ċE����Z����W��ʙ�ha�Аwg�_�`�noE�!��0������� �:~f��D ����1�q���Q��>Ou?W�uvl:Զ�x�W�m���Į���K��v�xa-�\L��d���O��l��͆���˽���C'}a�-�g�P#)�u�i��4錸�ؓN��6���xz{`,��.�3kݰ+Q7;�������h~�*kɪ�n: 0��?���>�3p�������m%� Fe#�()�qK���>���v��#���)�JgJ��=��g^�\
|
�HC�
�2����V������s�l�P�W=��](����#�'g96�!k��y��� �lT���*���Rɐ�:�y�J�`ri��h���Bp�
�G��o4�pu|ޣ���$%v�p��N��(�z����G��x�+2sP��8����a���=�v��p�˅x��A�Ȼ ���OK��rO�PfzgT)P;9���W\!�6/�T����,���P'���EC�a��K/��0d�5���M+����F�`������L���qbg
Xq�
cVǹ��@s��z7�%�b~����)s�����D�q8�KA�:�?�:��xtTO�{�R�;�A6�Z&��+�bț�B 6]�g�}Zh��;>��P�Q�ֆ�����#���r��H�U0���g�X����,<����.Z�y��h��el�o 	�&y���Hְ��ݱ��	T��/������^ �'�6J�x�ڧ����՛Jɡ>oZ]PtN�%���3C��R�3��^�S���nY[�С��鳐F��T}���u��-�-o�7f�5�����rʴ�/8>Cot��ee(�p����č\���� �LS�*��K��cQ'b�='��B�^�;C��sBo�Րz��y�b���	�nԬWp��t�E:��m����SW��z^m���[\^�67�B܋�Ŵ<���/�h���,��࿼�@
�����I%�O�H-�]O����:q�a`�
G��H�={	�k�`:N[T�6��j�S9!m�K���zH���)ϼ��g��s�
1\-��2`�k٨k��K��8�]}�+�t�2�b*DL �V8���V �^��]��mԋe�&M��q�%C�ь�;�˵%_#R��O�: ރ��-���Ƞr���@�ng�4!�&�)%5 �W?:;�O��fO/�E@��b,uyH��ohh��X ~��%e	���@���=��kF�);3�wh�aB0V7Q{a�aQ�BB���-9�(�Ԓ�X�(�-��R�u ;V�$�'���~�su--Ê1 ��Ҵ�|+��̹�m�/ո�a���[6JM��Q�x���<tB�U�C���w�HJ�Y圔	��Y�i�͑��>ws��>3�uB�Yѵ?�����(}��H/2c��^d��׊���ߋ�m�����d�$r�I��+��؄���YJh
.f��
�=�:�\��	[˥{9�\l�<|o�	,'9	p����|y1y�6 ��C!aX�\��`vz|!W�f�SO9�I�u�pf ��Ҍ�3g�D�Z4pH�9�}�����[|A��>skm�����d��b�6ٖ�%N�K�`x$@M>���FCu�Z��qGS�j|!��Z^�Hp��gg�h��a҄sٛ�6�tic~����3��	2�H���2�Y3�f:������r��^�N��k�*O1�Ycm'$ۆ����mCs�� {_��~J���Ld�0]��ik�ۿ�({L�"K�U���S�wӯ	�ٵ�+��Kx����QOɢ���B5�D>�Z۪�����l�rib�俒^6�_��[���򥾳'���羞Ƹ��[�x��:S�6���i
{Ė�
�2yfW�\	��i_�2��=�]5�rgȵ���_�3��M�Sa�� ��?�J��ݶ�M�m��Q8_��7/⨡�J�<�᫮���M���Ŕ%����ۨ/QB?V��'��U�>}�ا1*�Ac�$��y�����t�S^b1�oٌ�c��.5 L("��'O4��B�*�)7�,��ֻ�i� O�
�~�^�^,�!7 �Xj�|��F��C5v,���O<�_���~h�$�Ï�5�},>����Gr�l"H1jZ$ʕ��6��I����s+X�Λ��f�
��ɵ%s�9��c�����5���u�8�`w ��R�o���Q	ڲ�:��~p��9o�Ӗ >���\�E�
�K�:N�Ywү�2�����D��2�n~v�J�ѓ%T.)���u0���^ �X���5�6��ȓ�3���ˣK�j����ά�cEo��8���ǌUJ�hM�S��BF�Ӵ������0���U����M����/����h��4�{Z� ���0g�{�1 6�%O�/�������{*l5;��Y�7��D�D����5��X�<���MG]�q�Og��r��o�����͵�Bn����z���i!�[�'���q��{tst`oE'�.�	֦|q"��h�қ��Ĩ�t
I��,��K+(5���(RoYk�UҮ&"¢k(�x��2'H�y�̰Г�������/��p�^�t��<R_�b�P�g����s�g��nmm�4���V�K��X��֚g�-��Gs��BZ���'��u�]q��}`�T!�cV�.��lJ��h�=z�[%T6W��jX����x{mQI<�R��OG���.�ss�����<D��y����ޚI�͢�<���6�0���
������B����T�I�VM��'�
^u(�9���gX�<4
J��H�Y��b,y�p�ˋ�?���c�"8�Ĕ�!A��4�8�i�}$�]�n�$�R���nl1�Ck��լ�����1�sD/�*�_�4]vOc{�hN�mm�qu��D���>�-܋�&��Ȭ3<�wj�@�����=fa
J��/S��Ҥ��H�����l�ì��"zYwj��!,]��A�r���6DӜ ����48茇��[�<�5#�Y��W^_�eB��s"�wwG:(5����X ꃺ���ܩQk����x"l�)�1`S��ny����2��t���Q�=�!H�Ͳq�icm7�h�����K��L�]Пc�S+Q>�	�`�*���&:;"L���+�t�"��@�	ϵx��؎D���T�h�Ɉy����=��	�軓xUL�kaSJҔ�/��nv@(�U��q���q�W!�q�)��/�=$�h��ۄ$d�2�</��Ø��-͇J�G�xv(����5��la�P�^j�OSt������� ; ������Fcd4��tb+eiOл�I���&~Zhg���m٫ZIX5��SN�X˷��n���W�-C�{�5C_���O�ʊ��Ϛ��Z�.���\�)̱���@|��/9X�Fj�g�5t2�t�1�xkX�]�,@�aVik�����^g-��?+���HPs;�9
�4���!,wY8ّ&1M΅@Bh��2-�J�mʷ7�b#F/��,�Ibp��ǵ���u�.$���v����ax�R��j(3��)�yc���Q5�H~,2�(�L��	ta�i��ܕBݧș�k���̫R�YCFu7[��
ҷ�T��L�Ay���C��v����@�꬇��B��2#ڦE#T��E�H��:�
%�.u���}��z*ki[)�i|8ː;9���k-���vY�k|�B��3P2�f�����o���r*�F�=�43�W0��~OM��CB���t�/�}1�i�Y5;+`v������7�?}i�{���	Hb�U����ݓe[�3^��D5Uӱ��B�HE���R��"�x�f��L�>j�ƞ̞�p+�fO�5��;6���a{#>p�.3y����bdN�﫜!�R�Mi���(z�zz�tK2l�2�DA{��p���ݛ)������M6ɰ2�Fө׵�ӊJ�Ե��g�j�s�"���4�8 t�t�%5��$��nit.����VC_�����$�vݩ?�#���Sf5Exdp��$����6����||�Sx�F��6����E5��'?ﶁ�l�!o;��|�HSȀS>��K�Ja�X�c�(��|�����<>� ����U������}6����浄c+�X�m�HEQ�`E������c�D''�珎�����as�r��\���R�fC:��:� ^�J��mZ#�|�Ƞ���	�ub���)�^
#�a�s�H<6�r�������a�QS>t�O����$$K��5�X��|@O!M�P��K��7s��r��?+J!��e^i�G<Z?���Y9{
��A�h�	Bdb�;�QaVR�t�{���W>��^4k���Y
�h\ �%��j0��w������-F�c� ׾�N��e��4�r�I���I�s��0 �"�WA'v
)xz�v�3(۩�syp�`}�8dF�_֥%$um�:b�q�o�6�c�����C	ڔȨᔏW9��R�[R�T'�ɠe2��*�O5�E9�vQɛ9���H�	��zF�j����Q�]��>A��&��I-�C?b��s���8� r��!q�#��$��A
��?
3�o?�k�\�W�DSAT�?�.����r.n#�_�c0�λ��Ћ�Ll�{t�%1�P<[/X-����
¢�>�P�����L~�{Wa��0����Wd�Z�,K2N���%j�
m����S����	��͓޵�?Lŷ���B �|�^���CF��:�����j�,�zTitE?�{H�}�E�-4c�I��C�O~N��/Q|<]��_:6�/�p7?àر8�㑶��]�R����:��-:�>�g�F�����ڣ��n�
�� ��]�t����y>�#�6�ސ����m�>�W��w�V/�Eq�Ff�҉�О��۬yYQ�� ч粽�bKh��Y�A�#�����e�/�d���������p:G%�=����+�H��	��m~�	o��F��\���{�_�,)O9��:�Q���Z!�9C�6���/���AQú��O�����Çqݹ��Jy�Ł��1����L����R���Wh�	qw�*|d��	L�h`���Yxܷ�Ƶ�Q������gݴ�0W�\,[|j73�������:��alB���:"p�RՋr�p�f�Qth�ҵ�*����{���5�w��e@%)�����Yj[�R�6pZ�4��{W�}�gJ&�Qn�88j*�Ju�	���߸
����n�x�"o}�=������B�}*�g�������l�2����_��1���I����p��H|w ��|g���˞]��	�*����^��w&f^����t�ųv5��:
��)�@��Ԅ%&�En���'f�A�F�����3������PrT$¹������^M���JZ�ފ���.�s����� $�)&���ӻ~����pB2��V�P�J���䏂J��_��en�:��"�՘�º�����)��' ������1��zm2���K�9,�+n�X�i���Өxj�x���O�Fr�`~�o0f�=�s�n��û`FͮGe�+�n�{�h#I"<&�x����T]�v&��	�nik���A?�o{/
�=n��.��q�j�Ƭ6RR_1V�#	�AY(�*In���J��t�%ir��Z �D!>B�F9@���4)�D��'�ڡ+X;Y��<��X��+z�+�wm�Xʿ,������X
iՆR�^K�H׉�k�Za׆�dC����I�Y�G���t�"���0QП�!b��e*��_J�z��%��Q��C9 �-Ӏ�.'<�Bv\�C ���@]7���5(i�^ى8fU׼-d��˦W�+O�e��K7TƱy�%���q�P�d �AԞFjB�3Xb���c�d/JR)>e�ܻ�Ӯq�j���XC�&�\����6��ׁ����)c"}ͧ�]Z�O$��f��y!�޽e���!jq�QaL�Z�z6p����,ܲ��ԃ��o�J�����Zヨ�؛��ᚮx�_J]�"4,�5��w)�ms3Z�5��~s���	��H.$>>�����ww��=��E���'Q��\�j$�3�9�t_u�TN���֖]*�CYn�"X��x�4��W�;"I��l� �H�C6�d��_��ɒg���8�4��@�a���#G5;��)���a�w�0�!��
����v��&"&��2+�Q��F�X�9���\��@v�:U��I���](!]��YO)�V�ti_���Puc�.U�o�h�
@R�$�C��Ԥ�s��e#ʪ��)�ȵ!�ƴ���|�JH9�������E��� ��oR�\Hq
��6�X����5��C���`�ȫ�|t`LѬ$����������6^tX%C��+fց�sZ;+����l!�tϖ�j0͒'U}F&�U�h|���eH}���2���Χ���Ն�-!��,�8V���5|�����{�g��O�]�
u�C��s���B2e���3t��ؒ�V�:�@3/EJ�,�����5���m'Ji�;�Q��Ǉr�ף9$�v䄬������x��� ���u�\����B ����hO��t�C��[���Z�b|4�E�ž���k�����]xU`�S�m�U�p��`s��0t���N�i+��$0_��+��Ky.��->�5+E3P�+������L�����F�ˀY����m����o������$[{`�e����wmbm��y���hSM���y�g�P �W"�w�G[z`�bǓ*�x��<H܀O}77�d����a��o�U�{2A����!��}T�s��U]�W�MZv���� W��&����%��_��,ڡ"�������;��1�Z~(�?=���Y��������0)Ǘ�
�0]弉͋]�G�[ i�ș����4�&�{�F���:-�Ea�Y֣�9��+c~s-�{0}w��6��oC�{�,
�l�ZH�C7��k�ѷhUJ���d d-*Tv�&V�FK��/���n1�6>^F��m���Ylr���2���I��8��z��"�;Q�� C�F��Rj���J]a%U�}�ٛ�ƄL�:���[6�l�k
>�4��D�憉_lݴjM���{�+���#�S��nh*pR5�XӮ�}X�XC��T����W.���yBQ�)�eå�K� -��̋S�%�K$pL�BΗ�݌�������%�]��	2���(M;R6���axh0σfB�&�,ކ� V�q2'Xy=��+�Fi9�3Y\}2�g5�nrWć�n�Pt��<��2�a�,�I̶�����_�{5<]s�})0!$I8o����il���ٻ��!�!/��?�GZ���s��)O�r��(?��}��4��Yj9����(\yX�9O!S%�.���݆�&x������5�鄍i�g� ���b �PC�X�%M1mܛ� ��^�M_�Q�����
NJ~�:4�N���&Gb��/���.���\J�[v+r�*�( ��[$x!Aڜ5��/G���4�}V�����)�����Q|YԳa2�el^�����:1��'�����T+]��`��h�R��K~�����;��{JD�Ma�u��{;�����>�d�/B��{+fr��$&f�ރ���P%��DWl[�;dw����Ȕ�X_vW�l<��G�X�1�9)�M��nD��$�ƾm� ��<G,�-�&�f���G�2W��{o?p�ܲl�t��:3r䬄ӧ�`� <8��@r壿!�Y0��c�^��Gm|���#�'b��L^f3Uߟ��y�RmL�l�9��Oo��3�S��M���>q�=B�W!\ �2�7Uz��0{�[��|A��>��w��j |��\����0U�� ����*=�D��{Ph(���i=i=�����Jۃ=����yԋx���x�F�B���I*7C{l�����r����4�<�ڛ�� ����l���$�P�'*�r��He��i�P��J�mWs>*��^{������k�^�5�]��+432���h<�Y�Zf�^El�R�I;��9ޙx�N�ӓ��bwGz&�[(�YB�'J�0nIY�0!ڬT:d'm��o�lmZ���(e����z*� 岗�Vm�2��5{�>�j�k)��A���2��6��jS���\EñL����3�t��q�mG�8�� XYn�+;�	Bt���������߬p���}��
<Y_���^���\�M�wq���k<���w[B�z�(˦�	��Oǀ�(,G` La�3v��]��苝���
h�e���xXil��S]`�14�4ޕjT�)���C�Xk�6?�ƺE����a�(9��ޠ�ޥym��,�l߁�j�Dǟ��֟����DZ.�io�
z��²�D4r���Y��.�?f�0��p��L����Ph4,�V5�3J:��S�������)������)2�P�SA����� J]�-��8���iAa�O13]��¨<k���x+ړz��o�x0��"��S��'���֦��I��"�9���l����9�i}}х6W����,qf�k( ����/D�1�Lt&�7%ڸ�ę	On_�(�rMT����VN���Z/㸞?��?I3�lrw��tm4�	f�l�<չ,3F ���Βuݼ�,��nM���b��Z$��wP��$��]�g~�$|�yb}���dqX����֨�-�:���������R�gg��;-��p�P#ú����X��#w`�H[�߁�"*�D�gTCW���u��[�f�i����Ls��L�n*'��^7aGnU������w��$�y�b��e&J���,XZ�uyB��Ѻy�T� �Sز����O���\��}�9~j���Po{B{��Z$"�+D�J9���JJm�lW��e�����(h�|Y�\,/�p�����k�)ɮJ4	��!;0����[�`�To-e���j�$�&Hrd�C�/�J�-[����*��Iz�q5P�	�Ls�v�-s��!���C�F)XL0a��q{��3��^�
e���h��'�H��uԌ�7�Y�z�f�!o%IxR�s����wē\`�Kf��u�)*�~}~�ч5y��u����u��y���uy�1�A��̦Ǎ+6�و��4	���y���!R�d
Ak~����hj�:��]TfE7�m��℔�~�1ή����L�Vo�|�ox���.&����o����5��?BW�ndGc� 4;���I��\cK1��D9i��`��)k�E��0JC:+�M�$o�m�¥қ�0�?\�B�Yo��c�kX��sd��F�:����5�B{|�b�_oN�h��~��osvE[���y02C1��'YR�m�G8@!U�Zy�(A��XV� ��&Y�9zRYM0�x�˂2b41��	�6?�V�D�x�}�EPK���N��de��S��n�"�sW(�v+!��t��0�ܓ���v�C��v��V�t�9���q�R�Y���!�����G����̆r���e��C�ʬ�V8��l+AÇ�7֤�CO��}�aʢw��f�
�+�YH��v̇@�x
?�D�}�*���#��s u�I�9t yV�6R�CU�c~�R*���z������e�@$i�i��b���8�������R�X��'L $�ϻ��O���C�>���=��GD1��5d�E[ѣ���2�Z�Z$9OZ�y���fo�L�A�))>�.�l��16HsCa���π]47%��>=�n�o�j�43�U>�p�rz��9��?j�v�a�w��f�}��)u�ST�\��\�`x�2��k��z{��L&A췗n�hrF�t�P&%���v�[��"Ѕ��/�N��P>�j��:?�8�m:��&�����P8[��L�������'W���.O��&w�^`W�D;������8����%��M2�b#�O�½w���c�	�r�i�SiO���-��3f����w�,��}1��NoX�I��ѳ�q�8��T��xl�Uwv(|E���!bɊ� ��U�l!#�fn�Mr�EN�����%~�_�L?����.m��(���l����,5�LI'E�+)y�U_d��|�^��^٫�d�\��5޼����-�lH*[z p���oG�^��E��K��3\�>q1���w��>W?w8	4�![�,����mޔڍ���F�b��Q9�ˀO/qq&d����:���r5G�4�A3�r��9+G*�F>��l����@��^:����i��kz�9������e�;�7FԄg��,z_�3f'�	��m\��1�\-Ňm�)�e���C(��d�S7�m��Iܦ�.`�p�c]���.h�!~����,,ԯb5���5�X�i1̖2uA�s�f!�e[�����z�6ac���OV��������T����ѓ�!�$I�$32�ہS(��(��Kj��m]��p����\z6_~0uFݽ3��πn�yp(�[�z���D"����sI���Ѳ��;ni��|�:q��"V���'������}���O�VEb�J��904�au�ǵ�WAF��L����b�X.%\`�7���Vs~�%?!�e߷ij�Kt�]�W8�
�F����F&��=dq��Ap!�;��7�tf�-�vY`��@��6Jw��,˜Snb��_��Y�w�E���%�BJ!3*�V���G>J1'JWΓ*�3
� Ⱦ�
`CxO�_�s&�J�J�b/��6+ϱ��h{�M�'��#���D1�,��n%j�3v7xZ���[z��������"W[�y�~�$�m�rVy)�E��ƶNH�����$�.g[��"(�0y�1B�4͕��8�_/J��8�?n+�A����_��!0��� ���D۶=	ѡkPwXs��-+�����!6�U�{|��xɴݾ�KD�!4%�r��U�f�� c���*�������gX_Ȳ�o��N�|gh�ߣ0�ГC��A��^�T�����`'�^%(��J�X��9d�^���lx��ĜFR��-/���{9Ds�N���>Ä�Jr����k8
�u#�oR�g"y���� ��S	�~fD�����h;֡ұ��w��Nw�j�����-�Ŭ�V��$�~����b����Q���-����O�1�4�����(Y<"���U�M�S?��m�jY���zh�K��`P�v��g�����J��K�o٧tpx��s��Gg�>��_�A���B�:eE��3cf4�h�2�o�b2�0�
�]�������);�D�K���ML�X���5NZ� O�P�[�1 VK��H����a��
,����y*��t� ��a�r'�!X%��	�b�{YY{'_����(���jf��"^��섉��H�.��0@A5��_�I	����̩\t�J�\�%1o�ŅF �ӣP���0Uj���ݯp6év� ;���Y��8�!���3�3�r¹C�p{%����Y��?�KzA�J����z	^���I��D����4��a��z���j��v�X�j��{���z1; �K�G�l<�eshO���A�hWE�p����Λ3w�5� T�	ЂΜ�sL��C���'�l��}毟h�N�v�Z1��FsZ�C��l���ϵl��2�O"@��)l�o���Q*V��*��f���=j��B��&n����|�jXO+$� ҅-�~08<#��X�~oLJ��/�aK��l���ͯs|�K�@)��>�
c�{��.e�0��m��9�A�f��a��8`]���2ܻ��7��0΀k���E��	�X��qrJv�Y��y�����y�S�摽N\�iOl�^��)]�O߆�@�%��p�x�`�B�0$v_���ڬp��P/c�[�@�H�U�v��qZ��]�a�9�<��[�<&�g.GVa��VA*B�Q"٩oH�k> �at�ݭU���
�$=`:���W���]B}?��S1B:�}�q�����?y~Y��^&nAܭ�UWf���8�J�X8(���u3�X��P\�,�E��]M��w�.���)����HK�:7�
������7�*l_����ߘ%�7��OT��߲�����/�)Zf���$�Y�h'���t�P��u/���W!d�ҥ��=�+�*�9��z���E�w�q�1�0�g�/��o9!�
@�"t,����fV}F�r�!�~�/P3Z��f1=�ID>�h�Z��F*��Q��=����7_K键�
�U2�3�p��n���^]
KuW�0s�$�!Zn{�v[V�'Į��d���{���=���Ę����6.O�����<o��ի{��`�ӿ׻��e���?�Jc�H`��Q^�౅>yu��q�85�7<"�Q����GƊ�f�>u���Te����l���T��V�f��|b���W��X߻#ҥc�l��r]�3Y^�`K���(bl%P�IHd'v����ݕ�����N7΁��L���	��ҕS���$'5iL��S���+���/��D�PC�P��))C1���c`́�Q@B���Ⱦ�/31k���|��>�U$��*�G# ���i�l�.V�w�w7�-!c��a��/��NxӾS0��C��TwD)�C�Y�c)]]+SХ7Xx�R�W����&9�d �/Vї��y3n��-�3g"vH*X�\�����X��/�0��U�B��i`��{w*��F�v�O�җo+P��֠�T����t�ʡuƬn�`w4+��B�
�@dEq8��NZ�
L�d��nLG	���a! =I��Di���O"��9qin�� Բ�#%�TC1��e5��֦ ��T^����d��i�$���Ǐ��0�6���QFah��^S��BY�Ȳ}�H[lVɝ�ښ��jW<��i|ĩ���5��x��o�c���&�A��:�bi����~/	��J�&Zl�V��g�W�ʹ���Y�LRA���7�j��W��b3���6��E�U��bY��bwu-ՒO�韤?uP��;$��3�M9�l#��ܒ�-m��#��*y#���7��� ������1�f/FP�U&x?C"S�;�"����K���n��O�o�!����ȿm`�I�$����Z��񧟪~/�>d+-���2�_F���X�a���4m���M�JS-�9�������x?��l�46���N4�l1Z�I/J��z$ȶ������	R�k�:�Y���*���EG�.Q�Fם��2p��u��	��2����1��Z�������	e�nG�3�%�Ĭ���"��]�F����*'�ɉ81@��T��7*�đhp�oؽ�#���
��3��. O,�oD��^��^�������+O$-u;C��$KH���3x�|yA�&��t�]ћ��L����d�EO[	�V=Y�P�GȺa;����*�Ѳ�8��B�M�`D�}�Sx�+U93��;,	����-�r���O�J~�>����O�	?<Z*	��@�S�*\�b �҃Ky�s��aQ�q#��3�H$���'ʵM�tJ���8�Ƀ�Ƞ�>	4nc �9�^�4!^�k���Oc9/Ԟ\ҵ,�C�{Ѫ&~2>�E�%�� s<~��sW�x�[���\ئ0$�P�B�L8r��I���ő�!��Xz�d�wk̺G����w�����q�F���ߜ��F��Y&\sI��7��G��i��	��[j�STZ������_U�싆��
U[&}�����X	[/�S�י���@}U��\y W��\��U��w+���C�G�uj����_-���Z#_������6�b��N�M���wi���8��@V�Rg?�p�����y��!���I�<�\ɂ���f$f|!����%��z��ޙ|���S�����y+PxK5U�_�	��َ�o��o�#P赟�]�6��Ǌ�E����?jh`#4��4�<�Wug�/yI�}p�^)4��:����#�d��5���5|�ċ��������r��o����5F
�ȗ�x��8����fp�K�� �J�iߴ5�VP�6m��N��O���cmS�|�DM���p�E��̎��q���ӹJ�E�SY���u�F���4hƤ�x�Sd��(���8��Iyw*���Dǜ��-)~o���ev�9��%�����̀�9"IFX'F`[��>�
��`�0���Vh��D9������]
�
����a�6���{�L�ʳҪI�Rq&f�El��怄Kb{s��U����ٞ��`v���Px咆�����JI�82L`����]7��wRuQ�k� �K�ܗe_�|�H|-�Z�� ���X���,'6����#"A4>�����3fa��еVb}�`/�>�}��{cn8���;ӳ��u��	ƭ�}�f;a�P��j�\��F��ƈ�ԈtjU4?B�v��t	v<C\X~f�o'�ڪ��p�ʻ�A�\�fgT9ǻ&d6z��=��`����8�P�PX�kU�_w�A�v��M�|��0&j��j���ʽ;"ǈ�8�d��1��6ٝ2���{���Lf�k��C�V$j�5g�<Mܨ3'��U�U��Ψ%�Fg��chs^6��Nb)RM:�����|uwaw���d�6��6�vg'�[�@?*1f����ns�40������q�H��5fJy��m�e��{ �u�r"��-�s�'/��JZj@v�t`I�`�3�2����V�{���p�|�l��C�[���K1��9-d���
�uB"-���g������7��zs��CM���Z�5����@���
)��N�u2��w[�ࠒ�G��W�К7�o�qv߹r��1�9��������)�յ�xۉg|-�B�nN�*�}�:�_�.p�|Q+~d�f �tեQ��UV�c,��*2�Z�dH����@e�n���L� ���=0r�|��!��+��!rճ@�~�/h�L�윚�u����,���H�B�7�����\9������m�������?����6�2��pjF�\|�Sb&������ �I��|�Nuޒt����
&r�k.pܷ��7\")�0u��3��l��@���{�4J�K8ۡ�3)]g��!{%��%��;�傖��SJI�巳�D���N�����*�ͪu�I1�=������h�n�HD�y:wf�(�_�3����#�� �!�Hi��x� ��`lB�������̍-pșC���>�O�2�]	S�����L��>xM��}����?E.&9�V����[a5=X�`5��l�;L��o ���o���v�<�#��0�im`�d̯��s}0ވ'E{��E=O�E�I���`�\A�v���6�.C��;����X aُ�=y��8�Җ�$����9:i��pj�7+7��<6��k2D.�.Hb6(�����dq�;S�ߐZ*VF>R��nW{�<:$�;��y�a��(%̄jR�����Q��dI��*��]-��Fiu��)A�*���&��:-�g�<�Z��<��i����O�62��>�W���Qd�S?�H���Y�u�Tj3���7ùqf�� �&1�T� OÒ�	5���|������E��#g�ò�5+Ȋ�Ԉ��RHi��
H��Y�'aY������>�N�̆�0g�	d�$�W�n<Ұ��ʕ퓪�gO.���ua�E��t�2pg+.v�E1��m"\���Ғp��؟%,�.ܯ3V�q|q�k��r��<�t���4�����R90�9A2�m��̧�����+��č!8Y����v��:��x�`��{�έ穃�J�D�7����@��;�)�˧���6$u! �ǝ�_��Q�F;�D��Tf�g��-:��^��Ġ)���8���_7(��9�}�.��N�0

��2�ʚĊH�Zf0a)�9�F�>�%z4[|�8G��;t"s�nl��1�ˢ����ێ)�9,�;��
5|��}s7���%z�~)s�D��h�ϕ���!����T���C$��nlQ�0�����
K�vpQ�v4s�kz�#�Z��}%�[Ԫ��uH}�UUA>3piy@�w7�t'�rڎ�LUU2C6�%��j��l=z�E
�\M5�v��{�Cgl,ωK�8���Ϳ)���%Y霒�+�#c�l�����'i	���1� ��"�P�7d[���,����mF�4nǚ'�5��)Ʃ��B��Px'B5-��]�_ɱ�cg!pn�Ya��d��$]߳m�<�|�w'(pR�$�������Ä7/ܺ/����s�'���^˅�8�mά�%-V���	?,k=���v���v�;5�V�a5A��S1`�*<5�+���v�3�f�u8W�k@=K�D�[�˙�3�07��5!�z����������/�5h�7J�	⼼d�^t8�ڈ�HPT
��I_LRYI���qcL�k"� �s�j��R�C턙�q:���u��5��x�7�
?br�T�[ݠ�p�ynϣ�g���,8W��(/JVG #j�Zha��zG�Ԋ�*�*-����(�/?֢�$��C�90�$!�"���~�v��xt�/o�+aϱ�؜*J���v^!��\na
p���@r0������r�~C�Ճ]� wE��P
�����&Jj�Pob梇e��sv�Z���xi�?�@DѓhU��! �{rۺ��B��ir"/�����Ny��)�k�-��P?�k�f�I}�b&�$��x�=.m~{.`����ˎw�;���OgT�A��"!)N�ܸ1��*�*������zw��<9��,�l}0�b�]���U0��D���F���W�\��f6��|i;���Aa�J�nz�)�a�)�#C;�����z���ﱝ�4U�<e�b�]�D�e!�2��T�����}[;p{Q��,MX��k��n�`�*N��Q��Q���B�(��ګ�ٲ�xf�؎��R?Jt���v��Sh �=+�A�������SR���T������L:L�F�ؕ�*�@�a�,�#~l�Aq�A�S^���~շ�ZP����-�b����Ec5�W�Q�kPv�yx!i��d!^|/�Q���kI[�i�#�mU��5r�No�'��H�H��=�*�R��D��n��L<���CM�������J��3`@OO���'.k�Y�F>w��t��A�X�ie�|�B{E<j|���搠�=+cz7���EY��HvF���uf�f0��7@e���#�̜�z֣���#Z �!i~ț��D���cʫ�*7��z=Lu��b���������$��X��t\_���Ҿl
yW;ch�|��j\P�R��,`=�}�*���ٹ�BopeH�����!AX:��wq�nZ�/>t]W7t�����**��?󕆦ä�ѓR�+��@� p�Ȑ��hew[��O��SԸ��_��6eL� "r�z���e�s2>A�3��Dr\@�҅f����8������0�Ͳ����Ϣu��lE�dV�w����۴/�~�`N�e'��hpK�"�K�&��vDW0+���^��Jx���	�����z�qf �_��D�Y!��X�t�<�~��a;j��ߕb��{��o�܂�j�e[����9G��-z����~%0�c ���-B�?�Xm���C���Qo�m�s��/��xQ�&-L����+`+c��T��7�k�Qb �� Yn�'�t��P�.�݀�q{��d�$�3Ba����{_�_U�^��nU.���[�8t�gP2w���������� E��7������El�>�\f�Ty��ްb�mNwe�R[�*B����^�|��ջ�$�>x���󭗿��|��ʌ���E-�a�D���mGŴʱrB��}�m�i[LP��h��xq��}�&�z_i�q0��Yo�U�l �i�/ ǚ��(�$���n�c�T��rү �'9򀲮�lX�f���*ۥ��eA?��Ghʹ� :��l����Mb,�A�PAರ�R��ٕDVp��[_{�,��`�?�@�_��E�P.;�q�ߤ�=˦z��_ٚ2�gD�nu�nrb�6/�{ȵU�!��^g>^����k�T�<��:s�q���� q!� ���{����v |Q?���gۈ�xU��D뎍�vvlz�V�i����R(�TI���Aq@� S�w������+[������Ű~����d��&6?�._���>�4
*���ip����&��yn�ؚ�z�%��G�����Y������&���������͑��k��PK����p����S~_6]��0]�x�e��p�r��`��� '�����E�Z'@��Xy��]l��⭹�K�;Td;}Ó>�/@�dCAeD���H���Wd�M��^�۸'��!�R�F!���Ч��}�V����%�r�w�IS&�8�]up��\�{fpg��[��n��8�u�g�����Q|��OE��'�^��M�M�cDs-?�K�ӂ�y�2�6|�}ݯ��%�
Jq�CA U�x%�#��!)��p��1���3�Q���Z��oˎ(0��%&]�F5l��hTp��eMS���T���a�O=����D"9֚��DWH(�R�� ²�m����S���>M�Fݸm����mÂ�ԍ��I���A�����D�ܐ:핚��Ȏ��>x$g+г^p�O����H��`��؋;v4�F���3����ڵ� ���G�1瓡�+;��,����K�~����6���f(E$Ȧ�� ��ڎG�~Zx-'��)�����-�j�P*���C�#5X�Y6�u+��F�m�(O�՚T�*�zE�0�)���5_^�,�`P�	��-H��?�^�~����7�d]����,�˘��0`�V�/���R焻���_3�?��¹z�� �~�#�aZ1�}@[���$�W
 ~��v��֙{m9N����pO@�w��d~K����܁D�}F��$?���
ox(=�o�G�G�@���%�0�M��gR9�ٲ��.i�'k�&���*��2�'�᤻&/n��r��i�3��A Z1K7�~f̝����l������?�S���/B������B�1� j7�*-\�{������]��dX*(<I5w5l�D���&ζ*�#^�)P���DpC �Ga���;�6�*�Ù�*Z�C�J���!c2!�.�b�+��� z��r�_͢c���ba�N�kP�W}h��-s8����hB�&�~��P}"F�T�E�ړϴ�,���'$iX�
bδ��e@D��u���`�z�5���HJzo��+U��v{B�kg�b��.�\�3�>�*�!���W(�A��b�Cy�i���1Կg��Ā���.���%���e��]�c=�U��<_����I�o�zW��!�E�s�3�ꐷ\Ao�5�`�?V�5��Y�O���i�x#ϙd�`o+CאK��	:9ex:O T���>d�؛_|���rh�)��E�Pvj�m)��墘/ӀZ>�H����9'/���/�.�o}s���������EaK��������#�
x�Z{V���bc��|�s��s�V��쬉q��l��ɠC�D����b�� ��j����h��н���&Y���j_�5+b#W�Φ��b���x�����	y쭷~���4T��o 2_�rX�ľ�S��MI *��~��6A@>(�qkӰ�to�3���΄�RTJ�"F�H-�v��	�0'�#��[���L�S�� �PU}_��4���0�F��Čz*�����=Wv��|��g�����D]�	�Z )��)ʺa'8�ų�����6L<i��!��gL�r4�7Ƌ�3��Ӝh}Z��y���ρ�v���_W� ��1f�`Ŷ��tɋ�gL�5��ϝ/�^p�Rx�)d�����l9������㬥 $8��q���<
|F6����;G-��8�V�=���7g��I2A�0Y�[���nO��_=%\.�-��DߌM�l}�H�󁅐mލ���F���L�����H'Y�G��p�����n0;q.��p�2d���|KE��N��k��[��:����ȵ����h��+Ppb�'a��YhZٌ���\��BǕ�z��40]F~T��	�qp�o�~fs��<��[��o9�v�S'g�ff䵤�(�x��uN��j��`DM5���a��8����t��:�ۚ���u$�S/��6�2xJ��ƾ�|T�*��V��!�<�e�n@ �+���Ј�-��@��W*z����0]��,�x�'�9�LS�t$]��˅;��=N���ϱ��Y������nC����-"�_T�`����:ES�ѧ�S�k��2Q�؏ 9"�����̚�	�X��49���[Q�5�B���I�0ҧq�T�Y���{+;��	u���IR�IÄx�ԷN1�n���Pc�h��2���VZU�t��I9,�F��V���-\[P�)�N��ȡӥ��/5ւ ��Q��Ѧ=���`%�[�x��{����IH�Se��L^u�h'j�n�u�_)��&��l}���4R1����L��jb�����A�C-�8�4��0��s��G�-�"���S����`k]����/�.4X.z�1�`��Hd�:_F�
x=t�-�擻�*�~���,9_KUT������t���Ρ.����i��6B��	�!��M��$(;��+��wY�i�:�����e<�ze� ��x��w�'�J;�������=Gw��*1�����<G鵓���lm�F⥛3*���L�A�l|gr-J���#�/�G��O�����֯��)����F�I�a�/�B�"؇:�F�T�ION}= E�ymݓF�p2�����@�b@�4�3���!�y}A�f<���j�F�Wc����E�V9���� ��-���μ�DL`l0ȴ"��D�w�蛈 �M�|^�J��<�Sno�|%0,����]�['h"x���a#�@9�_�蹸�
\p�cg��E�9.(�O�Z�����`���DxY�M0�%���w��T3{( q��il�|L�2�l���BV_�*�FW��iLR6&�����eFB(L�#�y���.*,2v�[�/�o�����o��7���פ�=����f5�f����D�DSrU]��N�
�7a�~X<���nڻ�qW�`a1�jKOI�Pv��c�q�6|�;-l��]�V�z�x,=ϲ�6؅,�U������@�#X6�`yV��R�'m����;��#�2d������D3���8MGb<�>�@��'�@���@Xb�ф٣�`��aHYO���qTm�5�Q�s�_�i�O�]RA;�Ot��
s0�#T�n.U�ֻ�*��kN&	��%6T\r�\��jU���'�c�4��+�>��{�gG>�Ξ����
��J[𑭆lV�2N�|�n����R��(p��D�,���䳚u�"��41zx�hH��3h�(�0��RQ�?�0�eQ�.���� -v�Yf7_�pMRf����U��*,Y� 5�(j��C�9���.H�/����K�#�EӂeF� Dg�wNtN	�evb_T��g3�v��`�$�9~�ݜ���g��'eq#z����v�p���xYx�\�?���+�_,A��淚R�pJ�*&[��^ex(M����q��k�
�a�
�B?E�bj����u���v��Q圯�1N��VZ���" #���*5���ݞ5���P$o4T���"|kV�ȍ�Yz�h�쓞Bo6PvЧ�lV�D�i�zsd �8�	������t�X��s��ֳ0�̻����f3�ҧ�A\'�u�d��]�s�-�Ɨ&�B��ώ��x�G��������Gri	�x��I�u�Ʃ���;��Q��w9��5�t=�8Н���S�4�v�ٰ&k�9��FT�Cf���]ȉ�,�����$�0��O2�h��/jλ���F�EJdk��/aL���3y�+�8�;�8����l�?��2��p�NCm#��`ς%.�F}̀���Y�濶=R��ɫA�Xwᝡ�@�dǫ|�=I���T�Wj|�����{-�p�:��˱{;�\�@��j��k DV���D+М�N��� DN�[���z��Ʒ�y0�h8#�"���kw�'�J�ZX�f���`�M��Ӊ�TQ�c=�{>�Lu�l��é��{!xj����%�}%M��t���ͥf�K�4�0��A��U��}��0�r�R��N�.N������/�T�_ȹnO��w��o��.��#M��p2'Z+�pj��������w�V��1�ói����jb6���S��/��Lg�	��n	g�^b���b>|��zT�����*	Ry���,2QV�<=�:�
��������.<��c��
24�?-��7#_��^����`��q����1�g��O��v��g�|%�-�Q�m�k�_�<��,��'������q�7G�}/E�
�x���9|?Y鐔\S6M�dTb��zi����Ϳ1�2���t��'��Y{��7H��"F���2j����veƏ�e��dÖ'agF ��d}��U��#�ʋ�ܦ���:�\��	��7���&��M.�ջKrm��X��(��`n��w�'NC��S]�Li�L�T޽W�|�_��R���aְ��-_�0���|�#@hm9Mfՙ�O#��7��4`%���G͵d�g��<�F�S泆�iZK�x[pa���N�(a;��
�Q�����s'B6N��>���r"۠&��/�b�9
�r��֟��f��6��|��n_�8DN�
�o��շz�g��:�P-ݎ����L͗�<¢v��r�~ ����B3��@�1��"S�� ����h!�E��LǪ����Q6�,��"�T�q_PT�Ҙ:�b���ǼT:���2g�8P�D�&�3
��Nr�џ�N����	�{�����C]�xw��c��b�����{�Yb���o��z�7�v0�����&-���|�Z���ED�z���
ݏ�<u*ll�:��x�l.��̆&	1:�V�s�eX��Y�w0��NG����p
%��՘�'7�7�3=���t#��sg� U �oI�g,kkwT�a��L�c���Mj�z��.��T\B�A;����#X�����­�)����,�ᰕ �D��;$�[J/��h�j��4�kE�6Bپ��������Pͩ������s��3�n��'��68 /�tP-G��Ϭ[�}��_U�P�Z�wh�H�l)E�aq �
���Ph���c-��=v9NfC,�{��M2����>5��
-���X�D����h���&�̱1�i���X�4VL�ͥ�}P�V���}H�������\B�Wp��sC$#����h��S%Չ~�8F[<�˞������^��R���X�V9Ď��7�2W���D"r9�l�aZ����x�/i�9��m�G��%Z$]l�_����0`����ѸV�`��Sl}����Z�?#zwz(�Uv(�8��������ue[�J�����~����t����s���m�]�e-������l�<�>�h�~�?��/�/�:y'FMӶ�j�jq��Mdaw���:]}.ވrG�%i_���j��	��q~Ǩ��4݄��r���ҵ��4 sKwW��ZUax�&	nv,v��Z�O�^F�/W���
�9HyR;�a�I����?G#�:rbC�y\���8�?��Z��7�=c(p_k�XI�l�a��ȶ��H��-�jI����/�F�g�,Ǹva�¨��A��p|�޵)v��W��BQ�Q�+0��g$L���RU��$1��,Z�Ǣ%���$���u�7/�)�"��,OWT���4
<�>\�RV�h �6%V+��6��������Id��P���׺�͙KjjIZ�NH4�8����a�X���kS����M�}��Es�z\H�^R���խ������O���||2����q4���
/�+�q�L��A��S�V��8���\��1 �:[7�U�'6Lo��D�ݪ��~�s�(C���in��%�*��,���3���FU���HjA�f��S�
Z�}Ɠ�F�E邓�~~Gι_Swa�,��e�d��k"б��+8��K�+��f������� ?�H�>�����7�X![�����:������4c�1�#����|c�����s�gX�Hp�u�C�Y*�����[�����%7�g�i���~r�>n�kz�G_�i���~���x�^:�	����ܛ�pF0�#��v&-��K.��)J |!�!:H�߳�jDxTbQ<h	/Λ�?��9������Д^
����������Lg�?@�.	�[�pC[{עG�*At��
��O�U�̦�I��s*�|k����j </�|wU�#�ɳxM�G]��4ݪ��<�d3�~����Z͵"9�eX��jvEFNc�?yf��'��xnopj�U[�걕��z��NB�l_06�6��b��o+�Qe��	^��7.p�Lh�bL� ��+WNVe�8W�>�L�J���ߌ�K���#q(��^!����C��h-�4v,��2�2�pow�@�	�I\/��;�ȡ����@�P&P;���8Q�7X���?�}�l�����c��Q�N�'�6i��~���y��?,����+#IT/��\i*"P�l��|�".4�ͅ�r�ն^�ӂ�,�G�S|{�@�i��] Y�<Oӻ�#;��|��>c.6A�FT�96o�ߘ���C���Hy۶���Ew�'u�.�.%Uv�vxӌ���P#��[�B�y�#�RX���t��m�}p<u����MC�Go��\Σ����q�;4L�B�3!����z�q��.����eK���}�v;v�3��h�>>v���ݘ�g�hx?z#�"r��z>�=5Rے;�9>$8+Q%�ݠ8��vv뼲%�h��ǉX�Zq�������ݪ,럋d��d�׈�?[YE�Z�B�rK�?d�J�FE�1V�Iy���]��#h_����I5�J1`��3,ѧ��zw��T���+7s8���o�|	��-���a��4�g�s���!�c�MIb~]�Lt92�h�C��c�*�+�R�d8M�:�A�8�m����xv�sDܗ�{%pҢ�U�/��d�j�GJka\B7��sWz3e'�%ܢ,��-j��Y�"�A-6 3M�ߐn�O������0;_[�e�;�@x޻�齌h�K_���"H�u��v?����AK�5�Yw�UG	ze���[u�>���Hp�/���x򍷴��
 SW�e)�)�&)Bp{b�R#S��c_�e�Y4�svv�1��Z��D;�����:�~�P0O�з-&P"�R�v�vA���ܓi@�|������/��\(
�i0�*(�0ơ�vXdT$.�VK�Oa��_,�-p|��Jj�f�k����$Xv�9?������ҨP��_~9s��i��1�}pc����`��?M�����H铏��!�;|ZG�QL�I*��+"��lPS�$\��FO��Z	�aE&�%��SInm�F�v_n%_�w+D<�r��d��5���_~*�!���V_��> �X/�0 �ϖ���G�zȷ.���xC"�[�S��3��X�9��,}�py��,��yЊ{���<R�K( =�=,�ƽ�XaGAo�Q����fm$��9V�5��WϦd,�A9�8/~���%��/\o��oO���tn�G FX����)j�в*��P/	S��/F:���'��t�o?[�m5��E���b�����Fj�:�6.Y;O��up�N��="~���>O��j��)��tt)�QȽg4G��]�:ߑVD�O�p���Ͽ&=��_�V�s���Ir����o��Ɔ����Gd1�7iuk��sMd��8�a�N�������x����p�c�?a�f
��e��4j0�O<�]e�>]"�tl�=MC����Ң�7�p����e��ʘ��2�'u�r7����� P^��}�@�io�[ d�F	ʒ'���_@e�qضU�����Mi�xLا	��$G��b�*fX%�P��TC�E��SM���ܩ�zs/��������x{��v)|X��1�N�4m�cBXe��G�є�xI�Va@��<_�H�e4� BA ���/X�?2���^�5.1�v
�������s�?R��=������Gl�PM��c��Q����Ϗ� �B1b�6��SЬ��M�+����6�c^;���^Q~�0�����=���>�����V��9��
,�XW�������[4�bi�h5����W���ܱ��U�^鞘f[Cs׃h��SW�*}�w�X�5	6󰍗�q�^FQ��؂�m
7)�"ٽ�8)�>����5	��C���(��8�"kܙ<
@/d���1!l�1���8�SJֵ0�b��j�6T�,�Q|���<�r�B[��D0k��q��W��m�X0r�މx�����y/���b%N,�����o������|幙��6��;n��U����@��޷��T���js�[
���v���(��1�f�k�a��[�8k�ѝr5����w��OᕭP�9���U��(7�zǜz���S�_�����6�I��K���Z�%|!G�}��Xqx��t���3Z��/��_�6d�_�vAq��v�x#�X��*2��t�8�l<-�t�^�u�W��y'�2�t�� m�_�x���aY�����ō�@���m�XU��(R�#�	��?��^\�e?����@�M�]�q�K-)�]Ϗ�����n!#=#�w;~R�E ����k�u�����I�ut���n����W������1��+�G�s+���i9������%w��)���%d��{&���3'ﯗ0�e�ǹ�Hp��h 1��"��z.9�6d$��]������C�l)�d {[>�[��ۺas5�8�äy���DCHv5wu3���aL� ֆ�FUe�;Eh��
�)��;ڡe󱇞�D�|Q<�ُ}�%�j�kޚ/��x���RR���:�m�Q#OR寵�_��Nq�L�����@��P�NN��O�-��W���	�tq3~��Jk�Et�O��ZG�u�%�"�-�<���j�E�������4������u�]��7����-!5�9��w:3@��򓞌�0��:	~����!���y#(8�n+u��SL�7?,���_�����*?�	��!���YL�q騁�f��C'��DF�~	l�vY���nZIȓ�d0��##_�waۣ���r.�h!����s�a��i���~Qi*:y��Ix��� R(����0ѩ�h҅f�����Cˬ��M)WvX�&���¿U��`�hg�7����AR�>��IU���$C�1,t�o�	�[B̩nр�~~7y'x֣+�(?{���o�i{�	ƌӠ%�ǲ͵��D�tsmu�>GV^�������:����
n�_�s�2�/�pY��F����I,�0n��Y�\�0\���Umwl)�<l�3��YK>3��`�썃�bk�~�/��U[�z���Q|�z��"���}�!�x�.�+8�+?#�'��l�^���VJP7[:��w�-LR������&f3 �V�\��/�O�:s�im~/�s�GJ������R[L���Mc(�{��f0�&1�a&�Z5���QC��ND��N�?ӈ_�G.���
��q����JG�Ij��i��k��R���j��v;�l�O�[�1�p��+?��5K�(�T�T���Є<��F�_?qf�j{ԭ���3C�`�.�<�U�v��Cp�Z� #�/E+A�a��V(��Mo����o�C��GZi��˝f�#��8C��$�)ud��_����C�1ow��љ�>���:��盏g�� ]R�s׆Y���N��p�a^#��p=`D��
̜�[��ǆ���z�r�O?���%�5<�J��Tr$ݩ�-̭%f���VM\CJ��7�g(M7�j�R g��y���Y��)}5��IU��Q�8���Ԫ�9O�}ۺOD�VU����Ald��-26�̐lE�9��O�1��΢C0���3yFC�zS�e����ŵ)��':9��W��#�Y���B�zױ50�}b��ma��b���,}���MU=�H���1���]U0��g!�q�1��:\a�`���c��t麟�e����b���ђ�#^f)B�ia�,Tt�-��C!�(S����vt�ϩYSQ�#�_�O5�]T
�F�dTZ��+]ҝ���&ѻ�������W�sv��a�LiA�%�8�c�(�re�p�U�s?��-��2���ԏRc�R �D/꘳X?i���ebU\��*!����.�i]�ERe��J��gV��ۑ+TR3Z��F:o�Q;����z���'7��'ۻ"iӭ왻�V�+�T�Zb���|C*_4s��Ȇ{��������^D7����"4����%-�Ѷ���$
q��K����O���R?mz�j>Q��Y۪�i+{�z�Ss��ʶ�������Ģ�.�6��c�&�Ra8�t'U"�m��K$�݌L�J=�g�jM`�G2��w�]j�l.˂����(k�J���ܾ!M�HeV~�wʊm���tmU���dU�I����Ѯ	��ҟ>.G�A�L82���;�����9�(�Z��o0䴜k�/s�ε���ê����S��<n{7��|sWy��8$�J���d�=��ѕ����寑��}o��3���?� �s�m�1,��u����=BE�-  �I=oqV _�.�މ� QA���R6���ด}���:�� U�s{�.�����$E*��$_����J�n�m�Pĭ{�����g�H�L�4#m�x .E���9 ����I؁����R�^���3���ϧ�����s���Ƕ���3~qH���S
�ML�W��@( �l]�\��C�c��=q�U'���ٻC%c��q�-Uv���S+ʟp��~���V�4�!�3�"�(&f*���߸���ڏ���\V>uޒ��wpA*��B�W�9�#�p�J��뚃*�T����3�Mr���!��p���P@D���9fy�� ��&�0t:w�F �D�����Fk/�1�!(�;�#1�/��̣N�7����ɘ[m��g8���!L��4,!�t�W�O^"?��Pq5y���.�C]������&9�������$����n>	Jdɍ�o<y�e��d�U���DS�&dd0o��;-���+������+х�{n�"�҉��Z5�\��f2���'�}
"�I���85)�ϨHoq��W������[��T~�ޓ����_<Kt���Fc���;6�s �;a���&eQ��"�k9���UOw��C�Ή��E��RȻ��uE�Q��BB{��Ik�'e���Y��"�D����oW�2��]�O���¶�}B�O`*(}�	\���[Քl�"A�ɔ.��AG��c��U[ٛ�ޚ�Sݶ4���o��/KG�7F_��D働T�g�~���FW���jJ�wGQ�1�	�k(Wh�3Lrs������4�f� ĕPw�I���N�'@K�|5܁�6�X�s�h-�Uyy{:�D�����q��b#��)����|��{�?��سpc�*��>��1�oY�%;���2"�����)V{��7��2����`��cX{�\fR�_�%��&=/}�L�G�����mi��sS��RTP:�W��	��B#u�����y�Ԏ��������d����i�"(�Oh*:�,�K7J���
�S<Ce��\u:��u&�P������
�y
��O`��x�7>��q�Z��0V���YT<!�=!˩�_�0K-K�>4�[����Ђ��x/V��r~�U�Ĝ��,�5j�z/An=5���['u��j�e�fհL�GP�r���TT�X��6�pe�?�X����<2į�QyTܦ��$���貒�����0��l�g�w/x$K� kl�.^�ew[�AZ1�������ōz֨)�_qx�Y��5�����nc]<`���k�?}��H��v�^,���	�2K,�Y���}��t�W�,�U?y��1�V��p��/J�0T�Ʃ���o.�+ѕT9�hېlP��MPt���;.��`+��@�*h���
ȬC�5��&j0�p��ƣ������/eB�w)�M�2�hV죘�@rF6C�kб�ە��(�r�j G�6���A�b����iL��,���iA]���]P�4��C��J�(�����ɘ��]��P퇊	hm>�{�X>}�5~�����H'^�D�^A�덙��F�'���E�]�xf�lP|!�ؼpj�k�>Ċ�-1�y+W��J�����#9SG9^>�rː�֬g�J�j5͗�B �Nw�����*,� �.Q��u�	-���1�tm+�����5����v�Q��� d�����z$�88R����f��d���a�$��|��xr�ٲܦt6��"���P)�8m%��ZV����Ňj�Х����+M¼ ���z��T�r�BEV��E^7�^�nwo�zMKr�\�E@�r����.����Gk6�j�k�����w��� Ya��9Z+��H!c��.��{�� ��a�L��d[%���-�L�[V# �A�z�.V;�wۦ�K�Hm}h�o�I]㘮E
��J�C��(�/�i�C���S�  �	vJK�y�3ݘ*WP�I(v��7<� ��{���@G�0�v�e����,�.��Q�N���+�u�B:����������#���_˭�C���������8��D<�U� �i��Hr*�.����9��Z> ����[E�)M\���;w���MPA�9+9W{ߵ��k$�&��-�KZ:~�+W���յ+���W
s�皒�Ǥq�d����i��ҫ޷5&�5�%T���1�]���A�\��60N��/G_uR�����~�XA�sq�|P�Ͷ����O[��WI)-��|�)F�͔��a69z��ĩ��xdF��%��y��O���2.��~�{c"�%FBT-��L}� ����v�Ia�ȑ��*N�'�BY��gً���ظ�W�܄���56ik/j���8i���<ko�4Ι�..H1��?�:��ж�G�M@�M?�Ⳳ3�#<]z�oU�}i)�r7�lO�x��>�tq�
�Ds���i�l齇�M �I� �|����[��y�v��gM�e�*���lS�Yc�����a��!����ks��r�����b��s�YO�7*��z9^P��J����~U�p�k��p{���~Z�jx#?�̗�/�Tqi�/�r$
q�m�.��s3��U�W>�F��~��9p�Q�����b0��ۼrw�2���s�� K��6J�O�4����)s)}�{�ڋR0f�F�9�Ȉ~��=	�'����|6>�|���%�׹����Y7���M�"�L�([W� .�{7&E�xI�I������#ʗz�Y��A�\���~�|�k��)%k��e��T[sL�+�է+>a���pj��kJ�"u��"L�Y�2�xdOy)���x��CF�Ikv(����:��b
p"5Ȑ�th�!�,��C�eպ�P��<˻�����!��a�O8��φq?eUn�Qhճ|�mz��ɏ��-d���-��*������u<Z���g�"�Bي����\�G�h!��ݱ��ҳ}J��JB&�b�R�d���ٓ�c�wV-�I�*���~��E(3?H������p�n8��:O�l�B��z��k�A�[yD�)�j�O�@8�J>B6��ܡQebД��jܔ`��;*�0��)	d3:gX*kYxg'��)�J�s���E'��l��݄���&�W�I?h9�Ye�K��\�M���6�;J:	/F��˓&_�����(q6|�;��Γ\�%nd�s��o;�n�BHR�Q]���z�ㇴ���(<8_�/������h�8�H��];H_��n;=���Z8��Ų,ö*s�ĻQ'��Rq�R�M�`3+^����f�'��%4Rwݙ�H���Gv"����|m\:����>�6�ژA�u���Ư Z+1��٬?��r+&�2]��L;v4ތ
R������^�Y���^���W-�pVe�ᴄ?(��;	,�_M��]l���J^+�28��_����$6�,0�jO�V��S�Z�����n�8��>����q���Aa�g�
�O5���g��O
/�=��َ���^��p?���]�b��i��D��ň��z1e�����K>��`@��sG���F�z���"jՇ�"���pFG�\?$0�j0��
�w��+�K*. �����t3�kD���J�����K$wG�ڷ]��y�GZ���� ��I�}��!�T��ؓnD^��o\���x�h.g��|���">F���}��� ���r��J�-��sZ᧖��)"f����1�?\���NL"W�p�9acD�GU�Y�]��^8P�\�����3�+n>�$W�x���u!a��Eņt�?�S(�cI���)ӫ�}+�~�~K�ٰv����wޞg�É0�hM��kvgI.�8�ɇ�é������W�A1]Ǫ�2�-x|r(1�2�+�dL{��^�q�}�@�j�_����������	�G�!ʰ�-z�F���*eB�^��/P8a# S�Y�K梂@����@�ɹ2*̌�}���6�V�`��W��xCk�����{aD�@�]S�lyV��I�M���@T͝���hn01���R�m/@Y8�%"u�&�X@���ݕxb���i]�8�ҥ��/E��a�����������^3�J�F���
��ʈ��r`�L�>Y<��z�;��o��j�����������1 �}G�A�v⎱z]l@?Qp�j b��6�iM�j�������;W����d�������4�����镧5�/��y�W�2,̻���{�l*�%���B[�Zç� �%��}�+���:��L�Ƅ�9�G��t[�`�ԯ6SGɖ�&v�n^xo)J���Ơ�ˏ�\>�Q��z��:�za�҃1UU��]�=qi&v��ʎT��� �B������0/�U��ȓ�H�2y#9t �ǽ7`���}��˳�S1z��/57T~.��&�b�b���`���s�p3�uz!����}~�o�nm*e}���R (y���Do}ܾ梯�\����3��y��C��a�e@Q_�$9/�@��3Ԇ���W��z�.�n3�R�x�e;o��:���xA=l�.�m�5L�d�U�� �xY��"Z��֚��I�47Di�l���Lx��r��f�eί�F{<���b�}��|��]Z�������t�)��8;�� �Q�V��ܯj*���+ãy��_agr�3g�����D�UB�wVPe�]�;{`��Z����1{�����p7��1�jM�s'?���"�ʀ-W�Ȫ��_��ձ�T�r�$���'������x\/s�����L�-��~�u����2��u��cS��ק7C�i�A6�;��j�T���L�#�|뻠�]����c��4Qt(	t��Z�����#�Z�)�d{���.**��*���_-}�Ƭ�5��Xt��[5XJ`̰��ɘ��j��Q�����t%�wL�_�X�`�o#
5�� ڃ�zX������1U�-��/{*T��1������BmP[��8x���	��h΃rW��gL�m����G�E�f+��p������T�Ha1Ux��UC�t�c�K�o1}4I�����mH��#y�� J0�Xq҆0�v�x[kt�pW��"���HE1�T��3�?��j��L��L9lXnQ�MnG�Q˱��2��ɣ��[�>
��B;�ȁ��A��\SιyÓjPl������������\�P�`�Xd���y�׳\l	/} 4��~�F�U=[G�g���+��\/]�Z]N������lQ[�C����l~0�M��M�ɟ�̚s̝P���**J�	��U����^	�`���>�:T�%t��w�(��bfPx�?i?�� �2��{(u���a�����'\X�q\��s*v�����R��68ܝ8�b���Q���m�,�}k�ej+0%���G����%�I d
U�,(z�_h�����w�W�t!�&J�7G��U����
Ol$�}tr�����έ�]�s���^KkGaf &}5�k�c)���nlYZ���������$��J�p\��(�	��<��O�HP�\�_RRa�o���Q�K���,\R�")/3��#%�r���WeL4c�1$:�b�dc�$U�(B:-Yh�ct�f��u.����8�P��ˡ���1�Զ!�x�E���@K6;�ѧ-9�7���+�-E jO~�d�R�Y�Z�:����(��8�A��i�.��:%��:u�s���g�`�ZDGGw���g#_"�X�����&ǜ$iH��Kad�����%�`hKʂ�r��}Ě��E'f�:�M�zŕ����)_{���:�]��<%-K:���-�Y5=�=�M�H�k��`�S��)q�|�\P�c��-n��)���3�រ{@��j���l"��3��� ��46:��a+ѯȚԻn��#@#Dda�n�rN���DE����w��p+��4By*� ���V�|+`zb1AA����5]
�hI�����	LBz�:q�n����z��7;�M�9��T`� c�X��C5����%O��Bw�[�FpK,��� �%\����~�^�cl�j
�aIa[\�o#�����?Y�>�M[�Џ��H��Yes[���-&6��R-ڂR�äQgU]����Id�Pq�'�SH?"=԰&��}��S\O3��se�\PC �*8��QC��U���6�!r1+ƍHٷ����W}:w�@"nT�>���@��U��������9�;�u]b��
Ո1�4�~��]L����>�*Xݜsa��3O���NV! ��3���51��L�3�`-Њn|����yW�	\�z.�{�=ˡ�k��ߌ u[����L0%�A���Jb
���z��ŉؿ��(���xB�����
&�1��φ�$1X�%�����sR��d��辗���e�����ҍ�,�4=��+ҚpX�`�d����W�t �3��,J�iY�I�y	r��˼M�婙�� �j86v������+D�W��8�r��K��W�J,[c�j��4���W��w��=CS��R����q�l��]&�@�bP�؎}yA�&x����ЬI��J��#�x�^�g�n9r��'N���w������4R����5��J70�o^�F7��iGq�[�V?Ԍ�:�߈�Z^̣K�h�N#'����m����j�i 	��U݃B�B{/�j��{!'/
.�"��/��ۘ'����Z`C�v��E��<���cK�r#�s6JQLg�s^�7�d�D�|�����ɋ�nU�MmO�%,��Z@���@�@}ܯ��j�KY��M#�P�y�,WK���ZI�H Ls��9��%uK��>_n(��T�W�
 M2�J�?��l�A�;b�59xh�Zx���sJo���'r9�K���W��Ix�HBמܷ�B�$GFfb�o�Kb�*�����\<���. �V*�T�z��c�,���r�������K$B�Lu&Zb*���ip�!��;�i�P�����6a�7ωdZ���OeY����NE�H�{2��0���]>��M�ѕ�~�w{��:� !h��Dٺ���B0����@���gPsi���t(~� �r^*7U`��1).>̧/�=I^H)1ʠ�*�T�_J")O��t-���2&�c�{K��W����wB �T��O��.J�!��E���I��X�G�S��5*�ͪeRuJ�;H�q8=��j+y��
�)�<Tm3�aF.�c��1�`7�:[@j@@���4z��Z*���܉@I)[�f�=�ZP ��W:�+}�@aw�Lꤎ%�ё��f���l�r&��;�|{�c(�w�!��XC�v��N�b*s�a��'T�ԽyW���H����ӊ)0�^>�H�v��/%A�*��p�^I^R��9���{��
�	HF����{�ii�l`I�Ni��w�V�f;���_]��`��}�:I�Ou]ү��ϟ���">1��Sz��p,�TB�-��fa �ї�j�?��d���5��t �'�bb��m^�x�bA�G]���;8QV�n~��H��|S�F��t�]6�B��پf�[N�J���b>��|n�6k��[N� V�O��O_�z'ﭡ�( ��h�G�U�ޘK�\��5D�G�y��;*�^�͔����*yт��`l����`*�ZY�I��$q}�I`��^֏�@���u/�ͅgQ�C`��0�Z�a6�0G)ّ�]�J�6��R�M�CH�5�f�R6j�፺U��4�Ѓ��\�SK�Y���#.�\{1ۯ�X�)�5ϕ�YE	?��~T�Qlsr�,��+!=�DE���X��̌,C�X�w&������u�ɹ	 v>�S~�Q2����uМ�<���;f�6B<�:M>�@�8�ΡAk!{�h�"�δ�2.�������s�o?�$ xϝ10�0U�Pn���x��Xk���d�7 ,�AG*IU��(�F���F�
z���-o��d\^��*��ރ�4⯝�6���2*�0b��yh�{���L,V<#&�n���j�iÕ��#$��v�Z|A��?�Ň�i�o�t�}��V��(��u3r����{D6sy�{�+��-�l䩺V	J���O����!�{�Y�/#2]����!)bDte^�wW?+^4���%)�����ygF�����#sB��ꞧ�����c�Wh�l���t5:��ȏ~B�]�_L�9c�z�3@6�/����,�v�6$5߄K��oW��]�{ ���i0��ԇ�8�M����1sa[C���T�J�&�� 5洐������;,�I�����%^�� 栖�ե�'O�o�i2
�J1�iһ���\Y��8�	�Խ܊Wf��%LI�nG�����_5��鼂�s��cV�/�Z�7V%{��za���(�!:���}�6o]8{���E�ʾ�0�Y��H�K�P���U��q��4�*�+���ؔ��{�;�ᔷ�WEZۗjُ[���>�ꬡ[+NN_�[M`,sz�x[�� �Qgc@__���F��c�w�7m�/�Z/1���Ts��Y��k╿q=DH�b�V���_�{ ɋ*X�TŔ����sߣ��k��kv�+)�	�v�F���5<��,fG����gmen%�+�3�'�4dEIo��en]X����9�p/�'~>���]���X���@�&y��w�j��� �4�TgF�i��*4�"%{1IE ߾z\0B~�U�:��V\��A	�(�|����<�i���kS�U��7�VS	�H��u��!��uL�x$�c��{�_�a:4ݟ���S��VOv���sp�%����{ �(s�J����)f4��U��Z�G_�$��-O]VA����')�_WO�ɢu����~_�w�.���Z�o�`�ǥ�o��X��48G�[��X~~	]L]����Z;����a�
E��dy�3�Ac���5����SX�@u�%��6p�1�by�K�Q;bـy�!�Po�3�S0��^�)���.�o�����7o}��G>��9��X a�hfe3|��-��ʻ0|b�!�u�G�,b1����Q:Z�[q=ϊ�ÙY��#�w�1ɻN�sl
��<r$O�w���)n���4�"4UP��j�%FU��t�,���vCT3ܴܲ9��9=�oz�lEǌ�|��X�S��"��~��z�o��R�)��o�w�r�ˉ�yj�¨)�� *zEM��kO���9n=�}�9�_75��Z�K6U޳=2�Ni,�2xl*n#1P�2dUu'���k�s%���=�.�D��g ��z-3�]pa�l,��#D]���Q�{�w<7�E��� �D���eMeAVYa����*|4OD��8E_����s��cޝGڭTp���%�ꓞ�~2_1�+��r�Tx]��E|��\�ц��}-�%�H�~&<9�+�&Q��I~��c*HDI�Vb�8���T�F3���S�$(d4����w�[�[d���?^=�g1�mn��`�!+�P�k;�@H���O� tX��}&�+�"Kq<s2 x��G}B(��,��XS2�'�\�t�T�b�*O[iP"�l��|{�_Dq�!4o������ ��K�ir�I3�?u~���΍t��4ب���mgsg;�Q�Y{�ϧ�a�����uj}��X�(}vF��Z�Ohy{�v����<��q0�b*�i����8b�F�|)M��M��p�8Yڢ�����B�9�}�����8�ړM~��uzX֤��k�!�*o�i���!���n%��L,q��BrĎ��{]�_N��B-~��;H۸����|��Y]W[F�#a��~�LА������U!6XPv�kh�%"���6��o�kFƣ�;�*2䕴Y�ϑ��B��E/�rZ�9�R�=m�U(�Rc��0�~<����� �C���k�[?*3K�pr�芳y���Ki ���4�l�Bv�Y}6��Dk7x��T6� ;(���4��Z?�do����_�Tqv�H��6AE܉4e�u~�F1γ��GČ�R��/��~	e}d+O	*�+?��u��7�'���>P��ij�����9ӻ�3�`�H���9�zqF��I�Ъ�";f4m��N��
����gy�'+#�ݏ���1"���g٩����$;�c����*(o���p����5Ũ��l����������3/�J�>�̿�6��2.c��I�|/?ǡfڜ�{zv���I����nn��zOo�fl?���x?��R��U83��X�BU,�Fe�����G�R$АTh[�x�z{����)����?�Ih�����s��	�R�#�o� =���i�ρ�����W{�O�fb��}i���{c�Yi�EI$���+]���&
��,*y_�sx�]b��|89kT�B	�b-�Ɉ�	
lЦ��
�L����^%Mԑ�
K��/PihM�&R��Jt���8�kC)6�!»�*G�;ιq7Rf)�_D��[�;|�]��H��(T�D�5&Hԅ?ip�������gЦ{ZO�=Vqa��PJcTB��~W�������֒S�Z�l��ssS꜊�ݰ���`��[+=�,�A��W���O��>���ИOp����\9���w���̒��1~Qulh��\ʻ����,9�aX�L���(�Q�j/��i����CXv]�z�B�JzM`^����i��C���1�a��cͱrv���'	��T+L�oa]�*�Hߘ1׿���s5�"���k�N���^]�h��1-�6��g�t��)=�0[P�.)�иd��b!
-gO�D���=q��Y���iSl.R�'��n7������y�P�;B��#n7)Ɲ"�n�����7(��>�[�B����
�.��i{�!?��uB�^pY���Onb��P8t[y�T�O�t�W��NS_YT��)��v�BM6�|�ɎG�D��~��C>-@KJ�����K�+�;�{�)zQ�g�H�EW��x�4)A�a�� �S)8��`����7(��<��Ձ?�`L+N��8ґTPu��6��٦�������:Z�-�e�D#)H����\�vV�5�4��O�e)k�1<�,.������'���
,��:7��ܢa�|��6E��6�ᅺ-/�F�[�K|�u�Qdi	k��R��lvG��ڨB�ߦ0�^��e����QQ`��%Ʀ8+>E�?о����`�b��ͶR,=H���]VX�ڵӺe����w�r#`F��p��h���T_L�90^��W��	��#U^�0����^�B�T��ָ��,�)k:*�|޷(��Ɔ�]Sf�y����|����=�|+�F��I�Y� J�����G-~��h����'�Q�|ʛ\�?�pn�4�w��g��k� cT<�kg���$�|�b���K�%�+F�J4�@�lcq�i�-j�e��_�:CO�/��*�����&���zAW�Km�;���l�a�SU%~��p^���\�����]���5�\���L'�=�Fp_KV
G
���f>�"�d6;}��[�5�%��)�@;zO�!R@�A�d��FI�@9�rz�UZ%@��7�3�'��~��:�'����k_��a�9�-���d����z�5�*N��|��̹��=~�����a�@o%IʓQk�Rҧ��&zy[Y�̮��o5��{C����uk�>h��@~/��h�.��as�
h�����]��sѾe��^�0&|Ma�h�@k�z��c������W������*b~ӈ�(�"^�V뀙�丈<O*���9sr�ʴ7 �(�"~jO��D��&=j?��EpA.@�s��Er(��6�[�K��ndtJ`4A�ld�l1y�~d,KV�х��־as�8�Pa�ދ �r(b����&W�Rl��4-ي��L��{M��r-�!9+����ȼzmW��%D��|f�h�U&TK�Cj��� �T^#ɥ3rX/a"M�Qt����Feߏ{�-A������,)R�L��:��@���$�/~��l�!�NqOx�ۯĩ}���U-A�����.�i���>F��MeU����j�|���Q~Fm(�/a��cIE�4��	��#
��p {�����9����p��������b"&8ZsT���z=��uj7�e��Ab6j|���rq���S�� ���	//�����d��(�ǽ����f}���v�u�\���gĩ�l�^vݎ�-;8oڢ����)�3|9�S���[�t�t�qR,M�ZpY��ɑ�.�s��c��_�i������A���Ί8�3��r�P㯿b�� �&�"&͵*n�>z	b��IGۺA{��w��Ub��<���s�d����/̄�8���$#��/���$��E���Q�Ɇ�	c�\+��H�a�@�����3d�g
����6��>0Ю�]����� �́���S��mx>ᇯ� f,�Yq�f)\_bIq�(�Ka���Kj�c��a@=����4��ɬq��(�E��H��+)��[l����Ά��Tf�N��$���"A[���g@�:�o,�'X���'/���ߑi�L�	d�v�8��I�`�[��#��%��|�f::�R�G���f�#��v/���I5Lt�Jy�v��50��F&�C�)��-�Po8ٷg�tU����}��aIP��8y<@�ц���Ϗ 
�6d�/�	z|b��3=`(�`_Y��yBB����73q�̂�M9�O2\h3�5
n�J
��ه��u��}=�+P�t~�5I�PN�/�ך��\� ��O�$��@��°4פ��lc[�(=1���D�$�[zym��UOBo�LI��C�1�mu�=9;�5n�a��A|�
��{:���%�+�!��z������M�U23^�]�HcJ� tz{/D�x�]@�Av�7�(W@�����C�&��j��֫1V�N ���K�`��ۉX��;��@T��O����I����Y�s7;���)~cfN.?�����il�@�^�~���JqƐ�R-��<�Y�ZRӉ�K�`XA2�v�K�I�Sm* vP�)9����c�E�'�T�49���'!gH������.L�LC;k��\�n���${!Q��;	�	� S��A���u�6E|�Ag>$��Yl�F��OQ3��K���N�?�=מ K���Yt j
�h���nF/q�+������hK�Բ��۞۾H�@#3�LR(
��Ï��,�~�4YI��MM~������;/Zc��d��5�魏s�i��~��PJ8ƅe|�H{�;պC���ǨFqD�Ի�K��3��N@��v�^ll|m!!j�g���Ր�����z/@�Ұ�H��y�|n��P%�&|��#罇$K��<�X���ؠ9~<�v<)�2E�q�U���Yx�*gIm��NR�'".�0x��������`�j@Mڈ����V��B��`Bp?�I�g��G���<�,�	����7Z�{Կ�D�Nl����ͱ�q�pC5ǘ��(Fi0N3[
ԑN�sN����'֯�B?���_Jn�m_��R�����e/m��C�s#����O<��<��� �v��wEfГ �,��?g؃�eݖ)��x�JE�n�ݰB���D��G��m��v-�*���ڹ�=`���2�J)��}�y80�}$�ܔ.�� ��텏�J<�p�� �|��h�B��,���8�I	�D3�.�I�MC��7(?�~+�m���g��q%�7�8<x�~��n��C�h���v���
rY�+�{���H1#�%������(���2L���o6q\�	�Q|\�j�������|<�(��`�;��l�]��6BK��)��2)i�(P�5ιt�4�0X�iF	N~��:-�������>)5�o��<V.0��4d��p�t�IP���(y���;���{���>O��W�6׷�x����dTa\����:V��I�cC	?���}�ͣ:���ޫ��/��7J��-���E$�{Z��H|������	��@Df�1Q3����
�rS��K�d��X����|d y��v�Q6*�u��X!|���x�nl���R�6B�1��ϑ�!�Q��}�H�����kV��!I)qʞ~G��+�qW��H�E��V�;��!�S1\8r0j�=5d*�b�D���
\�PtM*��������#.�m�S �z�vejdu���pl�G/����\d�2��纜�@�B�>�4��	�G���v�zsr?�j^�Ȼ�=�h���?Ir.��#�3poޖ��e6 ��h���O�քd�ސKe;�MX>?���̌;��L�6����8]tw�=2�b�5�L������O=$�nQ�f6r�V N�j~�z.׷"��M��/߿f�p=W,���]AN�E�1�}��!O^�:���_\��y�Y~�%J�����tVޢ�{��������
�9C�}�(�l�V�1���yX�{�I�5�4�O��1y��	�� �t.b\d��4u��B��
��t�l�I����-�]p˱�o��'���%�$�#��<أ}��wQ{�m:(�}�����w(�W��+ŸV7s���@-Zk>j�ޜʦ��O�	�	���m���o6�έ�+�D�K݉���~L/�Ø6��V�<�b�G�bgt��"�	v]tx���C��� P��WNv�C������PE:�(��9��9}��Rg�:Z���� ��SD��)[���:��s��Z�\8C/�+��g��ɪ�n�,7�����7SLn�(�s}Ii"'�o3�-\k�<���>�h��6E���a!���>r��N8st�Tƚ����@�n���Lv���8RP	�I�����j�4�v�m��?������G!�YB $c1��t��^����ݽ�U�ճo"�b"������C
qHKN�X���խ%���}�H;�ѹ�:���᮸�a"��ƒ�>a`l���ٖf�fc^캙�V �2X]�˴�%� #�hN��%��ߞѕ��f�Z������dS#��Kƺ��P���rp����,����xb�9i�Ȱ\T)�d��#+���R{�%g�1"6S(���gg����"Z[9�6��\o�&Ƃ����I�r���P4A���(�e�N=��u��:e�pЫn.�Ud�����W�� ��_�#HyZ�b(�#�����'z|���	��-�;�_�� ~�HA��+�S��(�3�� #�VX0���D�HU�o1D.�+��i������G�<s鳥gX�yRR�V�6������.u!� 8V �U`�$C	m5�(ܰd��-�6l�^y�Zd�8Ս�	�E���,w�k���s�Q�)A(�G����Jx�K���>�]�5آWm�*�ƛ��vb	#߽юA���$�~�&6uT}�����
C菻7x�g��ݶmB���w �ޢ�m���mm�;U�,�v.#��[�I������"8��j��\�FR�����5�"X� ��my�
9h��V�ޙv���)8sLan}�1y��#�4�_�Q�}��df���Bo�.<��_E�/G+�)�Z&$��������î�Ih�RS����o<����|Mp�6��".3�@[�
���9�4��4:����"0ۧ1\�+��w�m5�^<��<	/���b����f�BCŷ������������U���C�=;�����;熃����>u	��`������#.Gc���g��]���`��&���" co��]������u�~Y�O����s6���N|��R�Z �xA�N��l�����"�;�䧜��E��o^�%��#�\�xS��a��I�VK�Y�z��-1���9�<r��%�}ʞ�N{9a�)��D�@~fcf��N���&ͨ[~;������>���ʐ��!�g^q�u\ ]h@ �����l������0?����-x�Q�9�A������m�(���G�[�#�Y�/�Y��e�^��7�ݗ&�_&ƹ���fC���#HW�Ng	�(��؅�MVx�t��"2�v���R�x.X+ܶ��<���B?�̵kE�Q���ӍW*qd}0,F�@<�?��A�=�i���X"�2N^;<���3�b��<��I�Pm�R���_����9-�y��!��iV�%��w���]=��.Xz;d%��\��f��l�<(՗l�]�rc��W��
�܋��oc������%��H�v�Њ�1p+BA��1
>`��@B�$�c�lN���i| �W����)���b'3&����+�4�E���iAy s��������<�ˈ�2�Y�_-1Ƀ| ��_��id�^gI�"�ل��o���(Օ:�ʲ�Dg��5�F�攣�ñzK�-s� �ZI��}O�Z(��b�`c��
�(�ra��׀Q�}8�) �T��KT�s� �!vh=C7ϩo��Zu�Y6�3��#�p�M$	�'Z��DyO�n�ϟ]�(�$zj��M2� 8L\�6R�y�y~}/�I�0�A�����󕡬C�����|抭�%j2�-�3�˱������QF�ٟ����hwy/0]�F�[_{Z��(ď�mƃ?3�$�:z�-+�[=�=i���Px?Xa���(0�Hg1�
�� V��-�	��`���)|B�����:��X�de�Q��^�E�`]���ݸ�H>#> �q��N�[��B��^O��EiO������	$ϩ�L�Ua�n@X��N> q�9�Z?����C���t&�	��lH>a�T<~��2��f< ^G�����6p�r�nW����կ���?���S����]�Җ���o��Eo�Hɡ�Y��ಒ�ĔU{�H�Sd�-Pį+������ܧ�&��Ei�7�5��+��o��)�� #ը�L�Z� ��2kb��IS�����4�XO*�(Q�f�n��������G��$t}F�rf���d���F4\Q�Cy�!UZ%�Y�hLV�3A�����ߠs����5���'�˫�8�a�kN�B*U-&�8����2Nw}��;���3*V��<Mi�lB뽿`�s���̚[���/���J�� O��nt ���m���L�k�)�! c]�-D�5���1��^JA`����1x��9m�j�W�5���Wj8������猁l�7x����/�W��|(u{����5��L����Wpy�oU�[ ��1�Y0�i�?�/��Aҡ�&�P�ؕ�j�����K���C#b\�_ђ^q��Xv������.h�QO�șr.�����h�<0 �m錅��+7}Vj:N��W]�߂�@#j�pU���;���V�����q�ib�9�x)����/�Ce�a-�+ɖ�x/^�L ��%��ئ5[ߞڟѫ�"i������o���W( �A9�i�Fݸ�G[ĸ �����-�,F�]lnN q���j���:!��-	�~�B����#b�{�ǽ9���<vV�%�\�d�E_
���@�"��Y��q�~�Gʗ�T�(n;�Hy_�l�Ѯga�8�X�U"N��r�1+ֶ5��	�)m}|��'"�<�Q�����&��ɔV��i��*��t�,���vf��ۜ�H�ٺn�\�~.2T��X�	�z�^��l��*��_$�&�!�Nb��ݯ��=�H�G�׬�@��G�����͒
�/�	�j���Df���j�t�sڕZw J���U���܅2���_0��x�ӥpADo��I���E�3g�j�{�2#��~ŝ�x��v�����q��O���v��b�{ӱ�
Z]��_ͅ�c�;2Sx���ZZ6�z�E/��5}O����p�E��Xڅ��U� 2iO�пӺ|�H�;2���:\��#�]��b��Jk��:���M��<�ee�_���l<���8{�7��,��Ad��HP>��+����T�aA��;��I��)H�zI�4U
~)|�c������Ҡ[����{�j�<q\��m�3)<+���� ��	m5�E�6A�u�S�)d|���C�IyΖm�\E�Y���Q��S$�d2nY�D��[���&E&���H��gj��+o�~8r�&�S�^ˤ�ӛVT8YV%U��
ԫ��s��������yt|���!0G\�̹}O Z��o����X<�j�x8&�)�|���"�Ty�U F6�s0O�?w�GOZ���x��7D�P��������Ҭ�R���μgt�-ې�>)$4���wY�)bF��b3By������U��u�������>�*6��6_g.�}�s���]�� �,3��'դ������H&Q��3-4B��O#�L�-����f!U)��vW.�6�.Mǀ�!��VJ�B.�6���(�a��Qt5	������_���2 �3����!�]��gS��B[F�d��n�,$u]\��1�)jx_����}��z	p�(�k��W����Pg	�(Րy�҆c��.K)���.��&٘Uf��٨�v8 >���~-���T8������wn��HbM��n0VG��n�Ļ0�6uO=���2�aZZ`�鎬���~q��̷��:�������!��F����~*���KJ"SI)�P�P̪��	�F���,FU�eɊ=Q��k�c��|Fϛ���'p����*���o��|3��,Uv�D�g �Ԟ)β.f���*o���:l������"��>�(m[o�a�)�� sM�f��K�߯>|�\q/�!�����݆����|�wO	6'rV�9�s��}�Z:qG�o*=t�Tj��9_���b'8.��*E���	����I�����D}j	zj5~���F��p�ڼ������e˼/7��6����L�Y=H1z